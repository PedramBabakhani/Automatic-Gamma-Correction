----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:26:01 01/15/2016 
-- Design Name: 
-- Module Name:    gamma_correction - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity gamma_correction is
port(  input: in std_logic_vector(7 downto 0);
       nrst : in std_logic;
		 clk : in std_logic;
		 enable : in std_logic;
		 gamma: in std_logic_vector(7 downto 0);
       output : out std_logic_vector (7 downto 0)		 
		 );
end gamma_correction;

architecture Behavioral of gamma_correction is

type look_up_table is array (0 to 252, 0 to 255) of integer range 0 to 255;
signal lut: look_up_table :=  
((0,189,197,201,204,207,209,210,212,213,214,216,217,218,218,219,220,221,221,222,223,223,224,224,225,225,226,226,227,227,228,228,228,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,244,245,245,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),
(0,181,189,194,198,200,203,205,206,208,209,210,212,213,214,214,215,216,217,218,218,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,226,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,237,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,243,244,244,244,244,244,244,244,244,245,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),
(0,176,184,189,193,196,198,201,202,204,205,207,208,209,210,211,212,213,214,214,215,216,217,217,218,218,219,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,244,245,245,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255),
(0,171,180,186,189,192,195,197,199,201,202,204,205,206,207,208,209,210,211,212,213,213,214,215,215,216,217,217,218,218,219,220,220,220,221,221,222,222,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,244,245,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,255),
(0,168,177,182,186,189,192,194,196,198,200,201,202,204,205,206,207,208,209,210,210,211,212,213,213,214,215,215,216,217,217,218,218,219,219,220,220,221,221,221,222,222,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255),
(0,164,174,179,183,187,189,192,194,196,197,199,200,201,203,204,205,206,207,208,209,209,210,211,212,212,213,214,214,215,215,216,216,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255),
(0,161,171,177,181,184,187,189,192,193,195,197,198,199,201,202,203,204,205,206,207,208,208,209,210,211,211,212,213,213,214,214,215,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,223,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,232,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255),
(0,158,168,174,178,182,185,187,189,191,193,195,196,198,199,200,201,202,203,204,205,206,207,208,208,209,210,210,211,212,212,213,214,214,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255),
(0,156,166,172,176,180,183,185,187,189,191,193,194,196,197,198,199,201,202,203,203,204,205,206,207,208,208,209,210,210,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255),
(0,153,163,169,174,178,181,183,186,188,189,191,193,194,195,197,198,199,200,201,202,203,204,205,205,206,207,208,208,209,210,210,211,211,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255),
(0,151,161,167,172,176,179,181,184,186,188,189,191,192,194,195,196,197,198,200,201,201,202,203,204,205,206,206,207,208,208,209,210,210,211,211,212,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255),
(0,149,159,165,170,174,177,180,182,184,186,188,189,191,192,194,195,196,197,198,199,200,201,202,203,204,204,205,206,206,207,208,208,209,210,210,211,211,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255),
(0,146,157,163,168,172,175,178,180,183,184,186,188,189,191,192,193,195,196,197,198,199,200,201,201,202,203,204,205,205,206,207,207,208,209,209,210,210,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255),
(0,144,155,162,166,170,174,176,179,181,183,185,186,188,189,191,192,193,194,195,197,197,198,199,200,201,202,203,203,204,205,206,206,207,208,208,209,209,210,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,229,230,230,230,231,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255),
(0,142,153,160,165,169,172,175,177,179,181,183,185,187,188,189,191,192,193,194,195,196,197,198,199,200,201,202,202,203,204,205,205,206,207,207,208,208,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255),
(0,140,151,158,163,167,170,173,176,178,180,182,184,185,187,188,189,191,192,193,194,195,196,197,198,199,200,200,201,202,203,203,204,205,205,206,207,207,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255),
(0,139,150,156,161,165,169,172,174,177,179,181,182,184,185,187,188,189,191,192,193,194,195,196,197,198,199,199,200,201,202,202,203,204,204,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,223,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255),
(0,137,148,155,160,164,167,170,173,175,177,179,181,183,184,186,187,188,189,191,192,193,194,195,196,197,197,198,199,200,201,201,202,203,204,204,205,205,206,207,207,208,208,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255),
(0,135,146,153,158,162,166,169,171,174,176,178,180,181,183,184,186,187,188,189,191,192,193,194,195,195,196,197,198,199,200,200,201,202,203,203,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255),
(0,133,145,152,157,161,164,167,170,172,175,177,178,180,182,183,185,186,187,188,189,190,192,193,194,194,195,196,197,198,199,199,200,201,202,202,203,204,204,205,205,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255),
(0,132,143,150,155,159,163,166,169,171,173,175,177,179,180,182,183,185,186,187,188,189,190,191,192,193,194,195,196,197,198,198,199,200,201,201,202,203,203,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255),
(0,130,141,149,154,158,162,165,167,170,172,174,176,178,179,181,182,184,185,186,187,188,189,190,191,192,193,194,195,196,197,198,198,199,200,200,201,202,202,203,204,204,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255,255),
(0,128,140,147,152,157,160,163,166,169,171,173,175,176,178,180,181,182,184,185,186,187,188,189,190,191,192,193,194,195,196,197,197,198,199,200,200,201,202,202,203,204,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,127,138,146,151,155,159,162,165,167,170,172,173,175,177,178,180,181,183,184,185,186,187,188,189,190,191,192,193,194,195,196,196,197,198,199,199,200,201,201,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,125,137,144,150,154,158,161,164,166,168,170,172,174,176,177,179,180,182,183,184,185,186,187,188,189,190,191,192,193,194,195,196,196,197,198,199,199,200,201,201,202,203,203,204,204,205,205,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,124,135,143,148,153,156,159,162,165,167,169,171,173,175,176,178,179,180,182,183,184,185,186,187,188,189,190,191,192,193,194,195,195,196,197,198,198,199,200,200,201,202,202,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,122,134,141,147,151,155,158,161,164,166,168,170,172,174,175,177,178,179,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,195,196,197,198,198,199,200,200,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,121,133,140,146,150,154,157,160,162,165,167,169,171,172,174,176,177,178,180,181,182,183,184,185,187,188,188,189,190,191,192,193,194,194,195,196,197,197,198,199,199,200,201,201,202,203,203,204,204,205,205,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,119,131,139,144,149,152,156,159,161,164,166,168,170,171,173,175,176,177,179,180,181,182,183,185,186,187,188,188,189,190,191,192,193,194,194,195,196,197,197,198,199,199,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,118,130,137,143,147,151,155,157,160,162,165,167,169,170,172,173,175,176,178,179,180,181,183,184,185,186,187,188,189,189,190,191,192,193,194,194,195,196,196,197,198,199,199,200,200,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255,255),
(0,116,128,136,142,146,150,153,156,159,161,164,166,167,169,171,172,174,175,177,178,179,180,182,183,184,185,186,187,188,189,189,190,191,192,193,193,194,195,196,196,197,198,198,199,200,200,201,202,202,203,203,204,204,205,205,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,115,127,135,140,145,149,152,155,158,160,162,164,166,168,170,171,173,174,176,177,178,179,181,182,183,184,185,186,187,188,189,189,190,191,192,193,193,194,195,196,196,197,198,198,199,200,200,201,201,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,114,126,133,139,144,148,151,154,157,159,161,163,165,167,169,170,172,173,175,176,177,178,180,181,182,183,184,185,186,187,188,189,189,190,191,192,193,193,194,195,196,196,197,198,198,199,199,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,112,124,132,138,143,146,150,153,155,158,160,162,164,166,168,169,171,172,174,175,176,178,179,180,181,182,183,184,185,186,187,188,189,189,190,191,192,193,193,194,195,195,196,197,197,198,199,199,200,201,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,111,123,131,137,141,145,149,152,154,157,159,161,163,165,167,168,170,171,173,174,175,177,178,179,180,181,182,183,184,185,186,187,188,189,189,190,191,192,193,193,194,195,195,196,197,197,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,110,122,130,135,140,144,147,151,153,156,158,160,162,164,166,167,169,170,172,173,174,176,177,178,179,180,181,182,183,184,185,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,197,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,108,121,128,134,139,143,146,149,152,155,157,159,161,163,165,166,168,169,171,172,173,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,197,198,198,199,200,200,201,201,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,242,243,243,243,243,244,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,107,119,127,133,138,142,145,148,151,154,156,158,160,162,164,165,167,168,170,171,173,174,175,176,177,178,180,181,182,183,183,184,185,186,187,188,189,189,190,191,192,192,193,194,195,195,196,196,197,198,198,199,200,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,106,118,126,132,137,141,144,147,150,152,155,157,159,161,163,164,166,167,169,170,172,173,174,175,176,178,179,180,181,182,183,184,184,185,186,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,104,117,125,131,135,139,143,146,149,151,154,156,158,160,162,163,165,166,168,169,171,172,173,174,176,177,178,179,180,181,182,183,184,185,185,186,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255,255),
(0,103,116,123,129,134,138,142,145,148,150,153,155,157,159,161,162,164,166,167,168,170,171,172,174,175,176,177,178,179,180,181,182,183,184,185,185,186,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,242,242,242,242,242,243,243,243,243,243,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255,255),
(0,102,114,122,128,133,137,141,144,147,149,152,154,156,158,160,161,163,165,166,167,169,170,171,173,174,175,176,177,178,179,180,181,182,183,184,185,185,186,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,197,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,242,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255),
(0,101,113,121,127,132,136,140,143,146,148,151,153,155,157,159,160,162,164,165,167,168,169,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,197,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255),
(0,100,112,120,126,131,135,139,142,145,147,150,152,154,156,158,159,161,163,164,166,167,168,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255),
(0,98,111,119,125,130,134,137,141,144,146,149,151,153,155,157,158,160,162,163,165,166,167,169,170,171,172,173,175,176,177,178,179,180,180,181,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,194,195,195,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,232,233,233,233,233,234,234,234,234,235,235,235,235,236,236,236,237,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255),
(0,97,110,118,124,129,133,136,140,142,145,148,150,152,154,156,158,159,161,162,164,165,167,168,169,170,171,173,174,175,176,177,178,179,180,181,181,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,194,195,195,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255),
(0,96,108,116,123,127,132,135,138,141,144,147,149,151,153,155,157,158,160,161,163,164,166,167,168,169,171,172,173,174,175,176,177,178,179,180,181,182,182,183,184,185,186,186,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,245,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,254,255,255,255,255,255,255),
(0,95,107,115,121,126,131,134,137,140,143,145,148,150,152,154,156,157,159,160,162,163,165,166,167,169,170,171,172,173,174,175,176,177,178,179,180,181,182,182,183,184,185,186,186,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,94,106,114,120,125,129,133,136,139,142,144,147,149,151,153,155,156,158,160,161,162,164,165,166,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,183,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,224,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,246,246,246,246,246,247,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,92,105,113,119,124,128,132,135,138,141,143,146,148,150,152,154,155,157,159,160,162,163,164,166,167,168,169,170,171,172,173,175,175,176,177,178,179,180,181,182,183,183,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,245,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,91,104,112,118,123,127,131,134,137,140,142,145,147,149,151,153,154,156,158,159,161,162,163,165,166,167,168,169,171,172,173,174,175,176,177,178,178,179,180,181,182,183,183,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,246,246,246,246,246,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,90,103,111,117,122,126,130,133,136,139,141,144,146,148,150,152,153,155,157,158,160,161,162,164,165,166,167,169,170,171,172,173,174,175,176,177,178,179,179,180,181,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,236,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,248,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,89,102,110,116,121,125,129,132,135,138,140,143,145,147,149,151,153,154,156,157,159,160,162,163,164,165,167,168,169,170,171,172,173,174,175,176,177,178,179,180,180,181,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,234,235,235,235,235,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,246,247,247,247,247,248,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,88,100,109,115,120,124,128,131,134,137,139,142,144,146,148,150,152,153,155,156,158,159,161,162,163,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,180,181,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,234,235,235,235,235,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,250,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,87,99,107,114,119,123,127,130,133,136,138,141,143,145,147,149,151,152,154,155,157,158,160,161,162,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,181,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,246,247,247,247,247,248,248,248,248,248,249,249,249,249,250,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255),
(0,86,98,106,113,118,122,126,129,132,135,137,140,142,144,146,148,150,151,153,155,156,158,159,160,162,163,164,165,166,167,169,170,171,172,173,174,175,175,176,177,178,179,180,181,181,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,255,255,255,255,255,255),
(0,85,97,105,111,117,121,125,128,131,134,136,139,141,143,145,147,149,150,152,154,155,157,158,159,161,162,163,164,166,167,168,169,170,171,172,173,174,175,176,176,177,178,179,180,181,181,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,83,96,104,110,115,120,124,127,130,133,135,138,140,142,144,146,148,150,151,153,154,156,157,158,160,161,162,163,165,166,167,168,169,170,171,172,173,174,175,176,177,177,178,179,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,218,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,237,238,238,238,238,239,239,239,239,240,240,240,240,241,241,241,242,242,242,242,243,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,248,249,249,249,249,250,250,250,250,250,251,251,251,251,252,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,82,95,103,109,114,119,123,126,129,132,134,137,139,141,143,145,147,149,150,152,153,155,156,158,159,160,161,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,178,179,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,237,238,238,238,238,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,81,94,102,108,113,118,122,125,128,131,133,136,138,140,142,144,146,148,149,151,152,154,155,157,158,159,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,178,179,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,236,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,253,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,80,93,101,107,112,117,120,124,127,130,132,135,137,139,141,143,145,147,148,150,152,153,154,156,157,158,160,161,162,163,164,166,167,168,169,170,171,172,172,173,174,175,176,177,178,179,179,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,238,238,238,238,239,239,239,239,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,250,251,251,251,251,252,252,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,79,92,100,106,111,116,119,123,126,129,131,134,136,138,140,142,144,146,147,149,151,152,154,155,156,158,159,160,161,162,164,165,166,167,168,169,170,171,172,173,174,174,175,176,177,178,179,179,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,231,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,250,251,251,251,251,252,252,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,78,91,99,105,110,115,118,122,125,128,130,133,135,137,139,141,143,145,147,148,150,151,153,154,155,157,158,159,160,162,163,164,165,166,167,168,169,170,171,172,173,174,175,175,176,177,178,179,179,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,240,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,77,90,98,104,109,114,117,121,124,127,129,132,134,136,138,140,142,144,146,147,149,150,152,153,155,156,157,158,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,176,177,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,238,238,238,238,239,239,239,239,240,240,240,241,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255),
(0,76,88,97,103,108,112,116,120,123,126,128,131,133,135,137,139,141,143,145,146,148,149,151,152,154,155,156,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,176,177,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,236,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,240,241,241,241,241,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,253,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,75,87,96,102,107,111,115,119,122,125,127,130,132,134,136,138,140,142,144,145,147,149,150,151,153,154,155,157,158,159,160,161,162,164,165,166,167,168,169,170,170,171,172,173,174,175,176,177,177,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,226,227,227,228,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,240,241,241,241,242,242,242,242,243,243,243,243,244,244,244,244,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,74,86,95,101,106,110,114,118,121,124,126,129,131,133,136,137,139,141,143,145,146,148,149,151,152,153,155,156,157,158,159,161,162,163,164,165,166,167,168,169,170,171,172,172,173,174,175,176,177,177,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,229,230,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,241,241,241,241,242,242,242,243,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,73,85,94,100,105,109,113,117,120,123,125,128,130,132,135,137,138,140,142,144,145,147,148,150,151,152,154,155,156,157,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,173,174,175,176,177,177,178,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,240,241,241,241,242,242,242,242,243,243,243,243,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,72,84,92,99,104,108,112,116,119,122,124,127,129,131,134,136,137,139,141,143,144,146,147,149,150,151,153,154,155,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,173,174,175,176,177,178,178,179,180,181,181,182,183,183,184,185,186,186,187,187,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,241,241,241,241,242,242,242,242,243,243,243,244,244,244,244,245,245,245,245,246,246,246,246,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,71,83,91,98,103,107,111,115,118,121,123,126,128,131,133,135,137,138,140,142,143,145,146,148,149,151,152,153,154,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,174,175,176,177,178,178,179,180,181,181,182,183,183,184,185,186,186,187,187,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,223,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,234,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,240,240,240,240,241,241,241,242,242,242,242,243,243,243,243,244,244,244,245,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,70,82,90,97,102,106,110,114,117,120,122,125,127,130,132,134,136,137,139,141,142,144,146,147,148,150,151,152,154,155,156,157,158,159,161,162,163,164,165,166,167,168,168,169,170,171,172,173,174,174,175,176,177,178,178,179,180,181,181,182,183,183,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,241,241,241,241,242,242,242,242,243,243,243,244,244,244,244,245,245,245,245,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,69,81,89,96,101,105,109,113,116,119,121,124,126,129,131,133,135,136,138,140,142,143,145,146,147,149,150,151,153,154,155,156,157,159,160,161,162,163,164,165,166,167,168,169,169,170,171,172,173,174,175,175,176,177,178,178,179,180,181,181,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,239,240,240,240,241,241,241,242,242,242,242,243,243,243,243,244,244,244,245,245,245,245,246,246,246,246,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,68,80,88,95,100,104,108,112,115,118,120,123,125,128,130,132,134,136,137,139,141,142,144,145,147,148,149,151,152,153,154,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,170,171,172,173,174,175,175,176,177,178,179,179,180,181,181,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,226,227,227,227,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,240,241,241,241,242,242,242,242,243,243,243,244,244,244,244,245,245,245,246,246,246,246,247,247,247,247,248,248,248,248,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,67,79,87,94,99,103,107,111,114,117,119,122,124,127,129,131,133,135,136,138,140,141,143,144,146,147,148,150,151,152,153,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,171,172,173,174,175,176,176,177,178,179,179,180,181,181,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,239,240,240,240,241,241,241,241,242,242,242,243,243,243,243,244,244,244,245,245,245,245,246,246,246,247,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,66,78,86,93,98,102,106,110,113,116,119,121,123,126,128,130,132,134,135,137,139,140,142,143,145,146,148,149,150,151,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,172,173,174,175,176,176,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,237,238,238,238,239,239,239,240,240,240,240,241,241,241,242,242,242,243,243,243,243,244,244,244,244,245,245,245,246,246,246,246,247,247,247,248,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255),
(0,65,77,85,92,97,101,105,109,112,115,118,120,122,125,127,129,131,133,134,136,138,139,141,142,144,145,147,148,149,151,152,153,154,155,156,157,159,160,161,162,163,164,165,165,166,167,168,169,170,171,172,172,173,174,175,176,176,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,241,241,241,241,242,242,242,243,243,243,244,244,244,244,245,245,245,246,246,246,246,247,247,247,247,248,248,248,249,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,255,255,255,255,255),
(0,64,76,84,91,96,100,104,108,111,114,117,119,121,124,126,128,130,132,134,135,137,139,140,142,143,144,146,147,148,150,151,152,153,154,156,157,158,159,160,161,162,163,164,165,166,167,167,168,169,170,171,172,173,173,174,175,176,176,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,218,219,219,220,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,228,229,229,229,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,240,241,241,241,242,242,242,243,243,243,243,244,244,244,245,245,245,245,246,246,246,247,247,247,247,248,248,248,248,249,249,249,250,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,63,75,83,90,95,99,103,107,110,113,116,118,120,123,125,127,129,131,133,134,136,138,139,141,142,144,145,146,148,149,150,151,152,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,168,169,170,171,172,173,173,174,175,176,177,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,215,216,216,217,217,218,218,218,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,225,225,225,226,226,226,227,227,227,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,238,239,239,239,240,240,240,241,241,241,241,242,242,242,243,243,243,244,244,244,244,245,245,245,246,246,246,246,247,247,247,248,248,248,248,249,249,249,249,250,250,250,251,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,62,74,82,89,94,98,102,106,109,112,115,117,120,122,124,126,128,130,132,133,135,137,138,140,141,143,144,145,147,148,149,150,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,169,170,171,172,173,173,174,175,176,177,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,220,220,220,221,221,222,222,222,223,223,223,224,224,225,225,225,226,226,226,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,240,241,241,241,242,242,242,243,243,243,243,244,244,244,245,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,249,250,250,250,250,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,61,73,81,88,93,97,101,105,108,111,114,116,119,121,123,125,127,129,131,132,134,136,137,139,140,142,143,144,146,147,148,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,169,170,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,220,220,220,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,229,230,230,230,231,231,231,232,232,233,233,233,234,234,234,235,235,235,236,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,241,242,242,242,243,243,243,244,244,244,244,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,249,250,250,250,250,251,251,251,252,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,60,72,80,87,92,96,100,104,107,110,113,115,118,120,122,124,126,128,130,132,133,135,136,138,139,141,142,144,145,146,147,149,150,151,152,153,154,155,157,158,159,160,161,162,162,163,164,165,166,167,168,169,170,170,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,218,219,219,220,220,220,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,229,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,243,244,244,244,245,245,245,246,246,246,246,247,247,247,248,248,248,248,249,249,249,250,250,250,250,251,251,251,251,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,59,71,79,85,91,95,99,103,106,109,112,114,117,119,121,123,125,127,129,131,132,134,135,137,138,140,141,143,144,145,147,148,149,150,151,152,154,155,156,157,158,159,160,161,162,163,164,164,165,166,167,168,169,170,170,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,228,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,242,243,243,243,244,244,244,245,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,249,250,250,250,251,251,251,251,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,58,70,78,84,90,94,98,102,105,108,111,113,116,118,120,122,124,126,128,130,131,133,135,136,138,139,140,142,143,144,146,147,148,149,150,152,153,154,155,156,157,158,159,160,161,162,163,164,165,165,166,167,168,169,170,171,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,221,221,221,222,222,223,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,244,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,249,250,250,250,251,251,251,251,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255),
(0,58,69,77,83,89,93,97,101,104,107,110,112,115,117,119,121,123,125,127,129,130,132,134,135,137,138,140,141,142,144,145,146,147,148,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,166,167,168,169,170,171,171,172,173,174,175,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,221,222,222,223,223,223,224,224,225,225,225,226,226,226,227,227,228,228,228,229,229,229,230,230,230,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,246,247,247,247,248,248,248,248,249,249,249,250,250,250,251,251,251,251,252,252,252,252,253,253,253,254,254,254,254,255,255,255,255),
(0,57,68,76,82,88,92,96,100,103,106,109,111,114,116,118,120,122,124,126,128,129,131,133,134,136,137,139,140,141,143,144,145,146,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,167,168,169,170,171,171,172,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,223,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,230,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,245,246,246,246,247,247,247,248,248,248,248,249,249,249,250,250,250,250,251,251,251,252,252,252,252,253,253,253,254,254,254,254,255,255,255,255),
(0,56,67,75,82,87,91,95,99,102,105,108,110,113,115,117,119,121,123,125,127,129,130,132,133,135,136,138,139,140,142,143,144,146,147,148,149,150,151,152,153,154,156,157,158,158,159,160,161,162,163,164,165,166,167,167,168,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,220,221,221,222,222,222,223,223,224,224,224,225,225,225,226,226,227,227,227,228,228,229,229,229,230,230,230,231,231,231,232,232,232,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,250,250,250,250,251,251,251,252,252,252,252,253,253,253,254,254,254,254,255,255,255,255),
(0,55,66,74,81,86,90,94,98,101,104,107,109,112,114,116,118,120,122,124,126,128,129,131,132,134,135,137,138,140,141,142,143,145,146,147,148,149,150,152,153,154,155,156,157,158,159,160,161,161,162,163,164,165,166,167,168,168,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,218,218,218,219,219,220,220,220,221,221,222,222,222,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,229,229,229,230,230,230,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,246,247,247,247,248,248,248,249,249,249,249,250,250,250,251,251,251,252,252,252,252,253,253,253,254,254,254,254,255,255,255,255),
(0,54,65,73,80,85,89,93,97,100,103,106,108,111,113,115,117,119,121,123,125,127,128,130,131,133,134,136,137,139,140,141,143,144,145,146,147,148,150,151,152,153,154,155,156,157,158,159,160,161,162,162,163,164,165,166,167,168,168,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,218,219,219,220,220,220,221,221,222,222,223,223,223,224,224,224,225,225,226,226,226,227,227,228,228,228,229,229,229,230,230,231,231,231,232,232,232,233,233,233,234,234,234,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,248,249,249,249,250,250,250,251,251,251,251,252,252,252,253,253,253,254,254,254,254,255,255,255,255),
(0,53,65,72,79,84,88,92,96,99,102,105,107,110,112,114,116,118,120,122,124,126,127,129,131,132,134,135,136,138,139,140,142,143,144,145,146,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,163,164,165,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,218,219,219,220,220,221,221,221,222,222,223,223,223,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,230,230,230,231,231,231,232,232,232,233,233,234,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,251,252,252,252,253,253,253,253,254,254,254,255,255,255,255),
(0,52,64,71,78,83,87,91,95,98,101,104,106,109,111,113,115,117,119,121,123,125,126,128,130,131,133,134,135,137,138,139,141,142,143,144,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,164,165,166,167,168,169,169,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,221,222,222,223,223,223,224,224,225,225,225,226,226,227,227,227,228,228,229,229,229,230,230,230,231,231,232,232,232,233,233,233,234,234,234,235,235,235,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,255,255,255,255),
(0,51,63,70,77,82,86,90,94,97,100,103,105,108,110,112,114,116,118,120,122,124,125,127,129,130,132,133,135,136,137,139,140,141,142,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,165,166,167,168,169,169,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,224,224,224,225,225,226,226,226,227,227,227,228,228,229,229,229,230,230,231,231,231,232,232,232,233,233,233,234,234,235,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,255,255,255,255),
(0,50,62,69,76,81,85,89,93,96,99,102,104,107,109,111,113,115,117,119,121,123,124,126,128,129,131,132,134,135,136,138,139,140,141,143,144,145,146,147,148,149,150,152,153,154,155,156,156,157,158,159,160,161,162,163,164,165,165,166,167,168,169,169,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,224,224,224,225,225,226,226,226,227,227,228,228,228,229,229,230,230,230,231,231,231,232,232,233,233,233,234,234,234,235,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,255,255,255,255),
(0,50,61,69,75,80,84,88,92,95,98,101,103,106,108,110,112,114,116,118,120,122,124,125,127,128,130,131,133,134,135,137,138,139,141,142,143,144,145,146,147,149,150,151,152,153,154,155,156,157,158,158,159,160,161,162,163,164,165,165,166,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,220,221,221,222,222,222,223,223,224,224,225,225,225,226,226,227,227,227,228,228,228,229,229,230,230,230,231,231,232,232,232,233,233,233,234,234,234,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,49,60,68,74,79,83,87,91,94,97,100,102,105,107,109,111,113,115,117,119,121,123,124,126,127,129,130,132,133,135,136,137,138,140,141,142,143,144,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,160,161,162,163,164,165,166,166,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,223,224,224,225,225,225,226,226,227,227,227,228,228,229,229,229,230,230,231,231,231,232,232,232,233,233,234,234,234,235,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,48,59,67,73,78,82,86,90,93,96,99,101,104,106,108,110,112,114,116,118,120,122,123,125,126,128,129,131,132,134,135,136,138,139,140,141,142,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,161,162,163,164,165,166,166,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,217,217,218,218,218,219,219,220,220,221,221,221,222,222,223,223,223,224,224,225,225,226,226,226,227,227,228,228,228,229,229,230,230,230,231,231,231,232,232,233,233,233,234,234,234,235,235,236,236,236,237,237,237,238,238,238,239,239,239,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,47,58,66,72,77,81,85,89,92,95,98,100,103,105,107,109,112,113,115,117,119,121,122,124,125,127,128,130,131,133,134,135,137,138,139,140,141,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,161,162,163,164,165,166,166,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,218,218,218,219,219,220,220,221,221,221,222,222,223,223,224,224,224,225,225,226,226,226,227,227,228,228,228,229,229,230,230,230,231,231,232,232,232,233,233,233,234,234,235,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,240,241,241,241,242,242,242,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,46,57,65,71,76,80,84,88,91,94,97,99,102,104,106,108,111,112,114,116,118,120,121,123,125,126,128,129,130,132,133,134,136,137,138,139,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,162,163,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,222,223,223,224,224,225,225,225,226,226,227,227,227,228,228,229,229,229,230,230,231,231,231,232,232,232,233,233,234,234,234,235,235,236,236,236,237,237,237,238,238,238,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,45,56,64,70,75,79,83,87,90,93,96,98,101,103,105,107,110,112,113,115,117,119,120,122,124,125,127,128,129,131,132,133,135,136,137,138,140,141,142,143,144,145,146,147,148,150,151,152,152,153,154,155,156,157,158,159,160,161,162,162,163,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,223,224,224,225,225,225,226,226,227,227,227,228,228,229,229,230,230,230,231,231,231,232,232,233,233,233,234,234,235,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,240,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,45,55,63,69,74,78,82,86,89,92,95,97,100,102,104,106,109,111,112,114,116,118,119,121,123,124,126,127,128,130,131,133,134,135,136,138,139,140,141,142,143,144,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,161,162,163,163,164,165,166,167,167,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,197,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,226,227,227,228,228,228,229,229,230,230,230,231,231,232,232,232,233,233,234,234,234,235,235,235,236,236,237,237,237,238,238,238,239,239,240,240,240,241,241,241,242,242,242,243,243,243,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,44,54,62,68,73,77,81,85,88,91,94,96,99,101,103,105,108,110,111,113,115,117,118,120,122,123,125,126,128,129,130,132,133,134,135,137,138,139,140,141,142,144,145,146,147,148,149,150,151,152,153,154,155,156,156,157,158,159,160,161,162,163,163,164,165,166,167,167,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,221,221,221,222,222,223,223,224,224,224,225,225,226,226,227,227,227,228,228,229,229,229,230,230,231,231,231,232,232,233,233,233,234,234,234,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,240,241,241,242,242,242,243,243,243,244,244,244,245,245,245,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,43,54,61,67,72,76,80,84,87,90,93,95,98,100,102,105,107,109,110,112,114,116,117,119,121,122,124,125,127,128,129,131,132,133,135,136,137,138,139,140,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,157,158,159,160,161,162,163,163,164,165,166,167,167,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,204,205,206,206,207,207,208,208,209,209,210,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,218,219,219,220,220,221,221,222,222,222,223,223,224,224,225,225,225,226,226,227,227,227,228,228,229,229,230,230,230,231,231,232,232,232,233,233,233,234,234,235,235,235,236,236,237,237,237,238,238,238,239,239,240,240,240,241,241,241,242,242,243,243,243,244,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,42,53,60,66,71,75,79,83,86,89,92,94,97,99,101,104,106,108,109,111,113,115,117,118,120,121,123,124,126,127,128,130,131,132,134,135,136,137,138,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,158,159,160,161,162,163,163,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,226,227,227,228,228,228,229,229,230,230,230,231,231,232,232,232,233,233,234,234,234,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,241,241,241,242,242,242,243,243,243,244,244,245,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,252,252,252,253,253,253,254,254,254,255,255,255,255),
(0,41,52,59,65,70,74,78,82,85,88,91,93,96,98,100,103,105,107,108,110,112,114,116,117,119,120,122,123,125,126,127,129,130,131,133,134,135,136,137,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,158,159,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,226,227,227,228,228,229,229,229,230,230,231,231,231,232,232,233,233,233,234,234,235,235,235,236,236,237,237,237,238,238,238,239,239,240,240,240,241,241,242,242,242,243,243,243,244,244,244,245,245,246,246,246,247,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,255,255,255,255),
(0,40,51,58,64,69,73,77,81,84,87,90,92,95,97,99,102,104,106,107,109,111,113,115,116,118,119,121,122,124,125,127,128,129,130,132,133,134,135,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,159,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,215,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,224,224,224,225,225,226,226,227,227,227,228,228,229,229,230,230,230,231,231,232,232,232,233,233,234,234,234,235,235,236,236,236,237,237,238,238,238,239,239,239,240,240,241,241,241,242,242,242,243,243,244,244,244,245,245,245,246,246,246,247,247,248,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,40,50,57,63,68,72,76,80,83,86,89,91,94,96,98,100,103,105,106,108,110,112,114,115,117,118,120,121,123,124,126,127,128,130,131,132,133,134,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,159,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,216,217,217,218,218,219,219,220,220,221,221,221,222,222,223,223,224,224,225,225,225,226,226,227,227,228,228,228,229,229,230,230,231,231,231,232,232,233,233,233,234,234,235,235,235,236,236,237,237,237,238,238,239,239,239,240,240,240,241,241,242,242,242,243,243,243,244,244,245,245,245,246,246,246,247,247,247,248,248,249,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,39,49,56,62,67,71,75,79,82,85,88,90,93,95,97,99,102,104,105,107,109,111,113,114,116,117,119,120,122,123,125,126,127,129,130,131,132,134,135,136,137,138,139,140,141,143,144,145,146,147,148,149,150,151,151,152,153,154,155,156,157,158,159,159,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,226,227,227,228,228,229,229,229,230,230,231,231,232,232,232,233,233,234,234,234,235,235,236,236,236,237,237,238,238,238,239,239,240,240,240,241,241,241,242,242,243,243,243,244,244,244,245,245,246,246,246,247,247,247,248,248,248,249,249,250,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,38,48,55,61,66,70,74,78,81,84,87,89,92,94,96,98,101,103,104,106,108,110,112,113,115,116,118,119,121,122,124,125,126,128,129,130,131,133,134,135,136,137,138,139,141,142,143,144,145,146,147,148,149,150,151,152,152,153,154,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,223,223,224,224,224,225,225,226,226,227,227,227,228,228,229,229,230,230,230,231,231,232,232,233,233,233,234,234,235,235,235,236,236,237,237,237,238,238,239,239,239,240,240,241,241,241,242,242,242,243,243,244,244,244,245,245,245,246,246,247,247,247,248,248,248,249,249,249,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,37,47,55,60,65,69,73,77,80,83,86,88,91,93,95,97,100,102,103,105,107,109,111,112,114,115,117,118,120,121,123,124,125,127,128,129,130,132,133,134,135,136,137,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,153,154,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,196,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,224,224,225,225,225,226,226,227,227,228,228,228,229,229,230,230,231,231,231,232,232,233,233,234,234,234,235,235,236,236,236,237,237,238,238,238,239,239,240,240,240,241,241,242,242,242,243,243,243,244,244,245,245,245,246,246,246,247,247,248,248,248,249,249,249,250,250,251,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,37,47,54,59,64,68,72,76,79,82,85,87,90,92,94,96,99,101,102,104,106,108,110,111,113,114,116,117,119,120,122,123,124,126,127,128,130,131,132,133,134,135,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,154,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,221,222,222,223,223,224,224,225,225,226,226,226,227,227,228,228,229,229,229,230,230,231,231,232,232,232,233,233,234,234,235,235,235,236,236,237,237,237,238,238,239,239,239,240,240,241,241,241,242,242,243,243,243,244,244,244,245,245,246,246,246,247,247,248,248,248,249,249,249,250,250,250,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,36,46,53,58,63,67,71,75,78,81,84,86,89,91,93,95,98,100,101,103,105,107,109,110,112,113,115,116,118,119,121,122,123,125,126,127,129,130,131,132,133,134,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,154,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,208,209,209,210,211,211,212,212,213,213,214,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,227,227,227,228,228,229,229,230,230,231,231,231,232,232,233,233,233,234,234,235,235,236,236,236,237,237,238,238,238,239,239,240,240,240,241,241,242,242,242,243,243,244,244,244,245,245,246,246,246,247,247,247,248,248,249,249,249,250,250,250,251,251,252,252,252,253,253,253,254,254,254,255,255,255),
(0,35,45,52,57,62,66,70,74,77,80,83,85,88,90,92,94,97,99,100,102,104,106,108,109,111,112,114,115,117,118,120,121,122,124,125,126,128,129,130,131,132,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,200,201,202,202,203,203,204,204,205,205,206,206,207,207,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,224,225,225,226,226,227,227,228,228,229,229,229,230,230,231,231,232,232,232,233,233,234,234,235,235,235,236,236,237,237,237,238,238,239,239,239,240,240,241,241,241,242,242,243,243,243,244,244,245,245,245,246,246,247,247,247,248,248,248,249,249,250,250,250,251,251,251,252,252,253,253,253,254,254,254,255,255,255),
(0,34,44,51,57,61,65,69,73,76,79,82,84,87,89,91,93,95,97,99,101,103,105,107,108,110,111,113,114,116,117,119,120,121,123,124,125,127,128,129,130,131,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,220,221,221,222,222,223,223,224,224,225,225,226,226,226,227,227,228,228,229,229,230,230,230,231,231,232,232,233,233,233,234,234,235,235,236,236,236,237,237,238,238,238,239,239,240,240,241,241,241,242,242,243,243,243,244,244,245,245,245,246,246,246,247,247,248,248,248,249,249,250,250,250,251,251,251,252,252,253,253,253,254,254,254,255,255,255),
(0,34,43,50,56,60,65,68,72,75,78,81,83,86,88,90,92,94,96,98,100,102,104,106,107,109,110,112,113,115,116,118,119,121,122,123,124,126,127,128,129,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,205,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,222,223,223,224,224,225,225,226,226,227,227,228,228,228,229,229,230,230,231,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,237,238,238,239,239,240,240,240,241,241,242,242,242,243,243,244,244,244,245,245,246,246,246,247,247,248,248,248,249,249,249,250,250,251,251,251,252,252,253,253,253,254,254,254,255,255,255),
(0,33,42,49,55,59,64,67,71,74,77,80,82,85,87,89,91,93,95,97,99,101,103,105,106,108,109,111,112,114,115,117,118,120,121,122,123,125,126,127,128,130,131,132,133,134,135,136,137,138,139,140,141,143,143,144,145,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,224,225,225,226,226,227,227,228,228,229,229,229,230,230,231,231,232,232,233,233,233,234,234,235,235,236,236,236,237,237,238,238,239,239,239,240,240,241,241,241,242,242,243,243,243,244,244,245,245,245,246,246,247,247,247,248,248,249,249,249,250,250,251,251,251,252,252,252,253,253,254,254,254,255,255,255),
(0,32,42,48,54,58,63,66,70,73,76,79,81,84,86,88,90,92,94,96,98,100,102,104,105,107,108,110,111,113,114,116,117,119,120,121,122,124,125,126,127,129,130,131,132,133,134,135,136,137,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,161,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,199,200,201,201,202,202,203,203,204,204,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,226,227,227,228,228,229,229,230,230,231,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,238,238,238,239,239,240,240,240,241,241,242,242,243,243,243,244,244,245,245,245,246,246,247,247,247,248,248,249,249,249,250,250,251,251,251,252,252,252,253,253,254,254,254,255,255,255),
(0,31,41,47,53,58,62,65,69,72,75,78,80,83,85,87,89,91,93,95,97,99,101,103,104,106,107,109,110,112,113,115,116,118,119,120,121,123,124,125,126,128,129,130,131,132,133,134,135,137,138,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,211,212,212,213,214,214,215,215,216,216,217,217,218,218,219,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,228,229,229,230,230,231,231,232,232,233,233,233,234,234,235,235,236,236,236,237,237,238,238,239,239,239,240,240,241,241,242,242,242,243,243,244,244,244,245,245,246,246,246,247,247,248,248,248,249,249,250,250,250,251,251,252,252,252,253,253,254,254,254,255,255,255),
(0,31,40,47,52,57,61,64,68,71,74,77,79,82,84,86,88,90,92,94,96,98,100,101,103,105,106,108,109,111,112,114,115,117,118,119,120,122,123,124,125,127,128,129,130,131,132,133,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,200,200,201,201,202,202,203,203,204,205,205,206,206,207,207,208,208,209,209,210,210,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,230,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,238,238,238,239,239,240,240,241,241,241,242,242,243,243,244,244,244,245,245,246,246,246,247,247,248,248,248,249,249,250,250,250,251,251,252,252,252,253,253,254,254,254,255,255,255),
(0,30,39,46,51,56,60,63,67,70,73,76,78,81,83,85,87,89,91,93,95,97,99,100,102,104,105,107,108,110,111,113,114,116,117,118,119,121,122,123,124,126,127,128,129,130,131,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,195,196,197,197,198,198,199,200,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,208,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,226,227,227,228,228,229,229,230,230,231,231,232,232,232,233,233,234,234,235,235,236,236,236,237,237,238,238,239,239,240,240,240,241,241,242,242,243,243,243,244,244,245,245,245,246,246,247,247,248,248,248,249,249,250,250,250,251,251,252,252,252,253,253,254,254,254,255,255,255),
(0,29,38,45,50,55,59,62,66,69,72,74,77,80,82,84,86,88,90,92,94,96,98,99,101,103,104,106,107,109,110,112,113,115,116,117,118,120,121,122,123,125,126,127,128,129,130,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,192,193,194,194,195,196,196,197,197,198,198,199,200,200,201,201,202,202,203,204,204,205,205,206,206,207,207,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,229,230,230,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,238,238,238,239,239,240,240,241,241,242,242,242,243,243,244,244,245,245,245,246,246,247,247,247,248,248,249,249,249,250,250,251,251,252,252,252,253,253,254,254,254,255,255,255),
(0,29,38,44,49,54,58,61,65,68,71,73,76,78,81,83,85,87,89,91,93,95,97,98,100,102,103,105,106,108,109,111,112,114,115,116,117,119,120,121,122,124,125,126,127,128,129,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,198,199,200,200,201,201,202,202,203,204,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,219,219,220,220,221,221,222,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,232,233,233,234,234,235,235,236,236,237,237,237,238,238,239,239,240,240,241,241,241,242,242,243,243,244,244,244,245,245,246,246,247,247,247,248,248,249,249,249,250,250,251,251,251,252,252,253,253,253,254,254,255,255,255),
(0,28,37,43,48,53,57,61,64,67,70,72,75,77,80,82,84,86,88,90,92,94,96,97,99,101,102,104,105,107,108,110,111,112,114,115,116,118,119,120,122,123,124,125,126,127,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,212,213,213,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,238,238,239,239,239,240,240,241,241,242,242,243,243,243,244,244,245,245,246,246,246,247,247,248,248,249,249,249,250,250,251,251,251,252,252,253,253,253,254,254,255,255,255),
(0,27,36,42,48,52,56,60,63,66,69,71,74,76,79,81,83,85,87,89,91,93,95,96,98,100,101,103,104,106,107,109,110,111,113,114,115,117,118,119,120,122,123,124,125,126,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,188,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,207,207,208,208,209,209,210,210,211,211,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,231,232,232,233,233,234,234,235,235,236,236,237,237,237,238,238,239,239,240,240,241,241,242,242,242,243,243,244,244,245,245,245,246,246,247,247,248,248,248,249,249,250,250,251,251,251,252,252,253,253,253,254,254,255,255,255),
(0,27,35,41,47,51,55,59,62,65,68,70,73,75,78,80,82,84,86,88,90,92,94,95,97,99,100,102,103,105,106,108,109,110,112,113,114,116,117,118,119,121,122,123,124,125,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,182,183,184,184,185,186,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,201,202,203,203,204,204,205,205,206,207,207,208,208,209,209,210,210,211,212,212,213,213,214,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,238,238,239,239,240,240,240,241,241,242,242,243,243,244,244,244,245,245,246,246,247,247,248,248,248,249,249,250,250,250,251,251,252,252,253,253,253,254,254,255,255,255),
(0,26,34,41,46,50,54,58,61,64,67,69,72,74,77,79,81,83,85,87,89,91,92,94,96,98,99,101,102,104,105,107,108,109,111,112,113,115,116,117,118,120,121,122,123,124,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,202,202,203,203,204,204,205,206,206,207,207,208,208,209,209,210,211,211,212,212,213,213,214,214,215,215,216,216,217,217,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,238,239,239,240,240,241,241,242,242,243,243,243,244,244,245,245,246,246,247,247,247,248,248,249,249,250,250,250,251,251,252,252,253,253,253,254,254,255,255,255),
(0,25,34,40,45,49,53,57,60,63,66,68,71,73,76,78,80,82,84,86,88,90,91,93,95,96,98,100,101,103,104,106,107,108,110,111,112,114,115,116,117,119,120,121,122,123,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,163,164,165,166,167,167,168,169,170,170,171,172,172,173,174,175,175,176,177,177,178,179,180,180,181,182,182,183,184,184,185,186,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,202,202,203,203,204,204,205,206,206,207,207,208,208,209,210,210,211,211,212,212,213,213,214,214,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,242,243,243,244,244,245,245,246,246,246,247,247,248,248,249,249,250,250,250,251,251,252,252,253,253,253,254,254,255,255,255),
(0,25,33,39,44,48,52,56,59,62,65,67,70,72,75,77,79,81,83,85,87,89,90,92,94,95,97,99,100,102,103,105,106,107,109,110,111,113,114,115,116,118,119,120,121,122,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,155,155,156,157,158,159,159,160,161,162,163,163,164,165,166,167,167,168,169,170,170,171,172,172,173,174,175,175,176,177,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,197,198,199,199,200,200,201,202,202,203,203,204,205,205,206,206,207,207,208,209,209,210,210,211,211,212,212,213,213,214,215,215,216,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,240,241,241,242,242,243,243,244,244,245,245,245,246,246,247,247,248,248,249,249,249,250,250,251,251,252,252,252,253,253,254,254,255,255,255),
(0,24,32,38,43,47,51,55,58,61,64,66,69,71,74,76,78,80,82,84,86,88,89,91,93,94,96,98,99,101,102,103,105,106,108,109,110,112,113,114,115,117,118,119,120,121,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,163,164,165,166,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,177,178,179,179,180,181,182,182,183,184,184,185,186,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,198,198,199,199,200,200,201,202,202,203,203,204,205,205,206,206,207,207,208,209,209,210,210,211,211,212,212,213,214,214,215,215,216,216,217,217,218,218,219,219,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,244,245,245,246,246,247,247,248,248,248,249,249,250,250,251,251,252,252,252,253,253,254,254,255,255,255),
(0,23,31,37,42,47,50,54,57,60,63,65,68,70,73,75,77,79,81,83,85,87,88,90,92,93,95,96,98,99,101,102,104,105,107,108,109,111,112,113,114,116,117,118,119,120,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,163,164,165,166,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,177,178,179,179,180,181,181,182,183,184,184,185,186,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,198,198,199,199,200,201,201,202,202,203,203,204,205,205,206,206,207,208,208,209,209,210,210,211,211,212,213,213,214,214,215,215,216,216,217,217,218,219,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,242,243,243,244,244,245,245,246,246,247,247,248,248,248,249,249,250,250,251,251,252,252,252,253,253,254,254,255,255,255),
(0,23,31,37,41,46,49,53,56,59,62,64,67,69,72,74,76,78,80,82,84,85,87,89,91,92,94,95,97,98,100,101,103,104,106,107,108,110,111,112,113,115,116,117,118,119,120,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,163,164,165,166,166,167,168,169,169,170,171,172,172,173,174,174,175,176,177,177,178,179,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,198,198,199,199,200,201,201,202,202,203,204,204,205,205,206,206,207,208,208,209,209,210,210,211,212,212,213,213,214,214,215,215,216,217,217,218,218,219,219,220,220,221,221,222,222,223,223,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,246,247,247,248,248,249,249,250,250,251,251,251,252,252,253,253,254,254,255,255,255),
(0,22,30,36,41,45,49,52,55,58,61,63,66,68,71,73,75,77,79,81,83,84,86,88,90,91,93,94,96,97,99,100,102,103,104,106,107,108,110,111,112,114,115,116,117,118,119,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,154,154,155,156,157,158,158,159,160,161,162,162,163,164,165,166,166,167,168,169,169,170,171,172,172,173,174,174,175,176,177,177,178,179,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,194,195,196,196,197,198,198,199,199,200,201,201,202,202,203,204,204,205,205,206,207,207,208,208,209,209,210,211,211,212,212,213,213,214,214,215,216,216,217,217,218,218,219,219,220,220,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,245,246,246,247,247,248,248,249,249,250,250,251,251,251,252,252,253,253,254,254,255,255,255),
(0,22,29,35,40,44,48,51,54,57,60,62,65,67,69,72,74,76,78,80,82,83,85,87,88,90,92,93,95,96,98,99,101,102,103,105,106,107,109,110,111,112,114,115,116,117,118,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,158,159,160,161,162,162,163,164,165,165,166,167,168,169,169,170,171,171,172,173,174,174,175,176,177,177,178,179,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,199,200,201,201,202,202,203,204,204,205,205,206,207,207,208,208,209,210,210,211,211,212,212,213,213,214,215,215,216,216,217,217,218,218,219,220,220,221,221,222,222,223,223,224,224,225,225,226,226,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,21,29,34,39,43,47,50,53,56,59,61,64,66,68,71,73,75,77,79,80,82,84,86,87,89,91,92,94,95,97,98,100,101,102,104,105,106,108,109,110,111,113,114,115,116,117,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,158,159,160,161,162,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,179,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,200,200,201,201,202,203,203,204,204,205,206,206,207,207,208,208,209,210,210,211,211,212,212,213,214,214,215,215,216,216,217,218,218,219,219,220,220,221,221,222,222,223,224,224,225,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,20,28,33,38,42,46,49,52,55,58,60,63,65,67,70,72,74,76,78,79,81,83,85,86,88,90,91,93,94,96,97,98,100,101,103,104,105,107,108,109,110,112,113,114,115,116,117,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,153,153,154,155,156,157,157,158,159,160,161,161,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,179,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,200,200,201,201,202,203,203,204,204,205,206,206,207,207,208,209,209,210,210,211,211,212,213,213,214,214,215,215,216,217,217,218,218,219,219,220,220,221,222,222,223,223,224,224,225,225,226,226,227,227,228,228,229,230,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,20,27,33,37,41,45,48,51,54,57,59,62,64,66,69,71,73,75,76,78,80,82,84,85,87,88,90,92,93,95,96,97,99,100,102,103,104,105,107,108,109,110,112,113,114,115,116,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,152,153,154,155,156,157,157,158,159,160,161,161,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,176,177,178,179,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,196,197,198,198,199,200,200,201,201,202,203,203,204,204,205,206,206,207,207,208,209,209,210,210,211,212,212,213,213,214,214,215,216,216,217,217,218,218,219,220,220,221,221,222,222,223,223,224,224,225,226,226,227,227,228,228,229,229,230,230,231,231,232,232,233,233,234,234,235,235,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,19,26,32,36,40,44,47,50,53,56,58,61,63,65,68,70,72,74,75,77,79,81,82,84,86,87,89,90,92,93,95,96,98,99,100,102,103,104,106,107,108,109,111,112,113,114,115,116,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,145,146,147,148,149,150,151,152,152,153,154,155,156,157,157,158,159,160,161,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,173,174,175,176,176,177,178,178,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,198,199,200,200,201,202,202,203,203,204,205,205,206,206,207,208,208,209,209,210,211,211,212,212,213,213,214,215,215,216,216,217,217,218,219,219,220,220,221,221,222,222,223,224,224,225,225,226,226,227,227,228,228,229,229,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,19,26,31,36,40,43,46,49,52,55,57,60,62,64,66,69,71,72,74,76,78,80,81,83,85,86,88,89,91,92,94,95,97,98,99,101,102,103,105,106,107,108,110,111,112,113,114,115,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,144,145,146,147,148,149,150,151,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,198,199,200,200,201,202,202,203,203,204,205,205,206,206,207,208,208,209,209,210,211,211,212,212,213,214,214,215,215,216,216,217,218,218,219,219,220,220,221,222,222,223,223,224,224,225,225,226,226,227,228,228,229,229,230,230,231,231,232,232,233,233,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,18,25,30,35,39,42,45,48,51,54,56,59,61,63,65,67,69,71,73,75,77,79,80,82,84,85,87,88,90,91,93,94,96,97,98,100,101,102,103,105,106,107,108,110,111,112,113,114,115,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,144,145,146,147,148,149,150,151,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,178,179,180,181,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,198,199,200,200,201,202,202,203,203,204,205,205,206,207,207,208,208,209,210,210,211,211,212,213,213,214,214,215,215,216,217,217,218,218,219,219,220,221,221,222,222,223,223,224,225,225,226,226,227,227,228,228,229,229,230,231,231,232,232,233,233,234,234,235,235,236,236,237,237,238,238,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,18,24,30,34,38,41,45,47,50,53,55,58,60,62,64,66,68,70,72,74,76,78,79,81,82,84,86,87,89,90,92,93,94,96,97,98,100,101,102,104,105,106,107,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,163,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,199,199,200,200,201,202,202,203,204,204,205,205,206,207,207,208,208,209,210,210,211,211,212,213,213,214,214,215,216,216,217,217,218,218,219,220,220,221,221,222,222,223,224,224,225,225,226,226,227,228,228,229,229,230,230,231,231,232,232,233,233,234,235,235,236,236,237,237,238,238,239,239,240,240,241,241,242,242,243,243,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255,255),
(0,17,24,29,33,37,40,44,47,49,52,54,57,59,61,63,65,67,69,71,73,75,76,78,80,81,83,85,86,88,89,90,92,93,95,96,97,99,100,101,103,104,105,106,107,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,155,156,157,158,159,159,160,161,162,163,163,164,165,166,166,167,168,169,170,170,171,172,173,173,174,175,175,176,177,178,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,199,199,200,200,201,202,202,203,204,204,205,206,206,207,207,208,209,209,210,210,211,212,212,213,213,214,215,215,216,216,217,218,218,219,219,220,220,221,222,222,223,223,224,224,225,226,226,227,227,228,228,229,229,230,231,231,232,232,233,233,234,234,235,235,236,236,237,238,238,239,239,240,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,251,251,252,252,253,253,254,254,255,255,255),
(0,16,23,28,32,36,40,43,46,48,51,53,56,58,60,62,64,66,68,70,72,74,75,77,79,80,82,83,85,86,88,89,91,92,94,95,96,98,99,100,101,103,104,105,106,108,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,163,164,165,166,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,199,199,200,201,201,202,202,203,204,204,205,206,206,207,207,208,209,209,210,211,211,212,212,213,214,214,215,215,216,216,217,218,218,219,219,220,221,221,222,222,223,223,224,225,225,226,226,227,227,228,229,229,230,230,231,231,232,232,233,234,234,235,235,236,236,237,237,238,238,239,239,240,241,241,242,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,16,22,27,32,35,39,42,45,47,50,52,55,57,59,61,63,65,67,69,71,73,74,76,78,79,81,82,84,85,87,88,90,91,92,94,95,96,98,99,100,102,103,104,105,106,108,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,154,155,156,157,158,158,159,160,161,162,162,163,164,165,166,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,180,181,182,183,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,199,199,200,201,201,202,203,203,204,204,205,206,206,207,208,208,209,209,210,211,211,212,212,213,214,214,215,215,216,217,217,218,218,219,220,220,221,221,222,223,223,224,224,225,225,226,227,227,228,228,229,229,230,231,231,232,232,233,233,234,234,235,235,236,237,237,238,238,239,239,240,240,241,241,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,15,22,27,31,35,38,41,44,46,49,51,54,56,58,60,62,64,66,68,70,71,73,75,76,78,80,81,83,84,86,87,89,90,91,93,94,95,97,98,99,100,102,103,104,105,107,108,109,110,111,112,113,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,158,159,160,161,162,162,163,164,165,165,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,177,178,179,180,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,199,199,200,201,201,202,203,203,204,205,205,206,206,207,208,208,209,210,210,211,211,212,213,213,214,214,215,216,216,217,217,218,219,219,220,220,221,222,222,223,223,224,224,225,226,226,227,227,228,229,229,230,230,231,231,232,232,233,234,234,235,235,236,236,237,237,238,239,239,240,240,241,241,242,242,243,243,244,245,245,246,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,15,21,26,30,34,37,40,43,46,48,50,53,55,57,59,61,63,65,67,69,70,72,74,75,77,79,80,82,83,85,86,87,89,90,92,93,94,96,97,98,99,101,102,103,104,105,107,108,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,152,153,154,155,156,157,157,158,159,160,161,161,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,193,194,195,195,196,197,197,198,199,199,200,201,201,202,203,203,204,205,205,206,207,207,208,208,209,210,210,211,212,212,213,213,214,215,215,216,216,217,218,218,219,219,220,221,221,222,222,223,224,224,225,225,226,226,227,228,228,229,229,230,231,231,232,232,233,233,234,234,235,236,236,237,237,238,238,239,239,240,241,241,242,242,243,243,244,244,245,245,246,247,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,14,21,25,29,33,36,39,42,45,47,49,52,54,56,58,60,62,64,66,68,69,71,73,74,76,77,79,80,82,83,85,86,88,89,90,92,93,94,96,97,98,99,101,102,103,104,105,107,108,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,136,137,138,139,140,141,142,143,144,145,145,146,147,148,149,150,151,152,152,153,154,155,156,156,157,158,159,160,161,161,162,163,164,165,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,194,194,195,196,196,197,198,198,199,199,200,201,201,202,203,203,204,205,205,206,207,207,208,209,209,210,210,211,212,212,213,214,214,215,215,216,217,217,218,218,219,220,220,221,221,222,223,223,224,224,225,226,226,227,227,228,228,229,230,230,231,231,232,233,233,234,234,235,235,236,236,237,238,238,239,239,240,240,241,242,242,243,243,244,244,245,245,246,246,247,248,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,14,20,25,29,32,35,38,41,44,46,48,51,53,55,57,59,61,63,65,66,68,70,72,73,75,76,78,79,81,82,84,85,87,88,89,91,92,93,95,96,97,98,100,101,102,103,104,105,107,108,109,110,111,112,113,114,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,135,136,137,138,139,140,141,142,143,144,144,145,146,147,148,149,150,151,151,152,153,154,155,156,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,174,175,176,177,177,178,179,179,180,181,182,182,183,184,185,185,186,187,187,188,189,189,190,191,191,192,193,194,194,195,196,196,197,198,198,199,200,200,201,202,202,203,203,204,205,205,206,207,207,208,209,209,210,211,211,212,212,213,214,214,215,216,216,217,217,218,219,219,220,220,221,222,222,223,223,224,225,225,226,226,227,228,228,229,229,230,231,231,232,232,233,233,234,235,235,236,236,237,237,238,239,239,240,240,241,241,242,242,243,244,244,245,245,246,246,247,247,248,249,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,13,19,24,28,31,34,37,40,43,45,48,50,52,54,56,58,60,62,64,65,67,69,70,72,74,75,77,78,80,81,83,84,85,87,88,89,91,92,93,95,96,97,98,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,167,168,169,170,170,171,172,173,174,174,175,176,176,177,178,179,179,180,181,182,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,194,194,195,196,196,197,198,198,199,200,200,201,202,202,203,204,204,205,206,206,207,207,208,209,209,210,211,211,212,213,213,214,214,215,216,216,217,218,218,219,219,220,221,221,222,222,223,224,224,225,225,226,227,227,228,228,229,230,230,231,231,232,233,233,234,234,235,235,236,237,237,238,238,239,239,240,241,241,242,242,243,243,244,245,245,246,246,247,247,248,248,249,250,250,251,251,252,252,253,253,254,254,255,255),
(0,13,19,23,27,30,34,36,39,42,44,47,49,51,53,55,57,59,61,62,64,66,68,69,71,72,74,76,77,79,80,81,83,84,86,87,88,90,91,92,93,95,96,97,98,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,116,118,119,120,121,122,123,124,125,126,127,128,129,130,130,131,132,133,134,135,136,137,138,139,140,141,142,142,143,144,145,146,147,148,149,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,163,164,165,166,167,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,179,179,180,181,182,182,183,184,184,185,186,187,187,188,189,189,190,191,191,192,193,194,194,195,196,196,197,198,198,199,200,200,201,202,202,203,204,204,205,206,206,207,208,208,209,210,210,211,211,212,213,213,214,215,215,216,216,217,218,218,219,220,220,221,221,222,223,223,224,225,225,226,226,227,228,228,229,229,230,231,231,232,232,233,233,234,235,235,236,236,237,238,238,239,239,240,240,241,242,242,243,243,244,244,245,246,246,247,247,248,248,249,249,250,251,251,252,252,253,253,254,254,255,255),
(0,13,18,23,26,30,33,36,38,41,43,46,48,50,52,54,56,58,60,61,63,65,67,68,70,71,73,74,76,77,79,80,82,83,84,86,87,88,90,91,92,94,95,96,97,98,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,116,117,118,119,121,122,123,124,125,126,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,154,155,156,157,158,158,159,160,161,162,162,163,164,165,166,166,167,168,169,170,170,171,172,173,173,174,175,176,176,177,178,179,179,180,181,182,182,183,184,184,185,186,187,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,198,199,200,200,201,202,202,203,204,204,205,206,206,207,208,208,209,210,210,211,212,212,213,214,214,215,215,216,217,217,218,219,219,220,220,221,222,222,223,224,224,225,225,226,227,227,228,228,229,230,230,231,231,232,233,233,234,234,235,236,236,237,237,238,238,239,240,240,241,241,242,243,243,244,244,245,245,246,247,247,248,248,249,249,250,250,251,252,252,253,253,254,254,255,255),
(0,12,18,22,26,29,32,35,37,40,42,45,47,49,51,53,55,57,59,60,62,64,65,67,69,70,72,73,75,76,78,79,81,82,83,85,86,87,89,90,91,92,94,95,96,97,99,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,158,159,160,161,162,162,163,164,165,166,166,167,168,169,169,170,171,172,173,173,174,175,176,176,177,178,179,179,180,181,181,182,183,184,184,185,186,187,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,198,199,200,200,201,202,203,203,204,205,205,206,206,207,208,208,209,210,210,211,212,212,213,214,214,215,216,216,217,218,218,219,219,220,221,221,222,223,223,224,224,225,226,226,227,227,228,229,229,230,231,231,232,232,233,234,234,235,235,236,237,237,238,238,239,239,240,241,241,242,242,243,244,244,245,245,246,246,247,248,248,249,249,250,250,251,252,252,253,253,254,254,255,255),
(0,12,17,21,25,28,31,34,37,39,41,44,46,48,50,52,54,56,57,59,61,63,64,66,68,69,71,72,74,75,77,78,79,81,82,83,85,86,87,89,90,91,92,94,95,96,97,99,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,152,153,154,155,156,157,157,158,159,160,161,161,162,163,164,165,165,166,167,168,169,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,181,181,182,183,184,184,185,186,187,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,198,199,200,201,201,202,203,203,204,205,205,206,207,207,208,209,209,210,211,211,212,213,213,214,214,215,216,216,217,218,218,219,220,220,221,222,222,223,223,224,225,225,226,227,227,228,228,229,230,230,231,231,232,233,233,234,234,235,236,236,237,237,238,239,239,240,240,241,242,242,243,243,244,245,245,246,246,247,247,248,249,249,250,250,251,252,252,253,253,254,254,255,255),
(0,11,16,21,24,27,30,33,36,38,40,43,45,47,49,51,53,55,56,58,60,62,63,65,66,68,69,71,72,74,75,77,78,80,81,82,84,85,86,88,89,90,91,93,94,95,96,97,99,100,101,102,103,104,105,106,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,136,137,138,139,140,141,142,143,144,145,145,146,147,148,149,150,151,151,152,153,154,155,156,156,157,158,159,160,161,161,162,163,164,165,165,166,167,168,168,169,170,171,172,172,173,174,175,175,176,177,178,178,179,180,181,181,182,183,184,184,185,186,187,187,188,189,189,190,191,192,192,193,194,194,195,196,196,197,198,199,199,200,201,201,202,203,203,204,205,205,206,207,207,208,209,209,210,211,211,212,213,213,214,215,215,216,217,217,218,219,219,220,220,221,222,222,223,224,224,225,226,226,227,227,228,229,229,230,231,231,232,232,233,234,234,235,235,236,237,237,238,238,239,240,240,241,241,242,243,243,244,244,245,246,246,247,247,248,249,249,250,250,251,251,252,253,253,254,254,255,255),
(0,11,16,20,23,27,29,32,35,37,39,42,44,46,48,50,52,54,55,57,59,60,62,64,65,67,68,70,71,73,74,76,77,78,80,81,82,84,85,86,88,89,90,91,93,94,95,96,97,98,100,101,102,103,104,105,106,107,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,164,165,166,167,168,168,169,170,171,171,172,173,174,175,175,176,177,178,178,179,180,181,181,182,183,184,184,185,186,187,187,188,189,189,190,191,192,192,193,194,194,195,196,197,197,198,199,199,200,201,201,202,203,203,204,205,205,206,207,208,208,209,210,210,211,212,212,213,214,214,215,216,216,217,217,218,219,219,220,221,221,222,223,223,224,225,225,226,226,227,228,228,229,230,230,231,231,232,233,233,234,235,235,236,236,237,238,238,239,239,240,241,241,242,243,243,244,244,245,246,246,247,247,248,248,249,250,250,251,251,252,253,253,254,254,255,255),
(0,10,15,19,23,26,29,31,34,36,39,41,43,45,47,49,51,52,54,56,58,59,61,63,64,66,67,69,70,72,73,74,76,77,79,80,81,83,84,85,86,88,89,90,91,93,94,95,96,97,98,100,101,102,103,104,105,106,107,108,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,131,132,133,134,135,136,137,138,139,140,141,142,142,143,144,145,146,147,148,149,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,163,164,165,166,167,167,168,169,170,171,171,172,173,174,174,175,176,177,178,178,179,180,181,181,182,183,184,184,185,186,186,187,188,189,189,190,191,192,192,193,194,194,195,196,197,197,198,199,199,200,201,201,202,203,204,204,205,206,206,207,208,208,209,210,210,211,212,212,213,214,214,215,216,216,217,218,218,219,220,220,221,222,222,223,224,224,225,225,226,227,227,228,229,229,230,231,231,232,232,233,234,234,235,236,236,237,237,238,239,239,240,241,241,242,242,243,244,244,245,245,246,247,247,248,248,249,250,250,251,251,252,253,253,254,254,255,255),
(0,10,15,19,22,25,28,31,33,35,38,40,42,44,46,48,50,51,53,55,57,58,60,61,63,65,66,68,69,70,72,73,75,76,77,79,80,81,83,84,85,86,88,89,90,91,93,94,95,96,97,98,100,101,102,103,104,105,106,107,108,109,110,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,127,128,129,130,131,132,133,134,135,136,137,138,139,140,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,158,159,160,161,162,163,163,164,165,166,167,167,168,169,170,171,171,172,173,174,174,175,176,177,177,178,179,180,181,181,182,183,184,184,185,186,186,187,188,189,189,190,191,192,192,193,194,194,195,196,197,197,198,199,199,200,201,202,202,203,204,204,205,206,206,207,208,208,209,210,211,211,212,213,213,214,215,215,216,217,217,218,219,219,220,221,221,222,222,223,224,224,225,226,226,227,228,228,229,230,230,231,232,232,233,233,234,235,235,236,237,237,238,238,239,240,240,241,242,242,243,243,244,245,245,246,246,247,248,248,249,250,250,251,251,252,253,253,254,254,255,255),
(0,10,14,18,21,24,27,30,32,34,37,39,41,43,45,47,49,50,52,54,55,57,59,60,62,63,65,66,68,69,71,72,74,75,76,78,79,80,81,83,84,85,87,88,89,90,91,93,94,95,96,97,98,99,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,118,119,120,121,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,152,153,154,155,156,157,157,158,159,160,161,162,162,163,164,165,166,166,167,168,169,170,170,171,172,173,174,174,175,176,177,177,178,179,180,180,181,182,183,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,197,198,199,200,200,201,202,202,203,204,204,205,206,207,207,208,209,209,210,211,211,212,213,213,214,215,215,216,217,217,218,219,219,220,221,221,222,223,223,224,225,225,226,227,227,228,229,229,230,231,231,232,233,233,234,234,235,236,236,237,238,238,239,239,240,241,241,242,243,243,244,244,245,246,246,247,248,248,249,249,250,251,251,252,252,253,254,254,255,255),
(0,9,14,17,21,24,26,29,31,34,36,38,40,42,44,46,48,49,51,53,54,56,58,59,61,62,64,65,67,68,70,71,72,74,75,76,78,79,80,82,83,84,85,87,88,89,90,91,92,94,95,96,97,98,99,100,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,136,137,138,139,140,141,142,143,144,144,145,146,147,148,149,150,151,151,152,153,154,155,156,156,157,158,159,160,161,161,162,163,164,165,166,166,167,168,169,170,170,171,172,173,173,174,175,176,177,177,178,179,180,180,181,182,183,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,197,198,199,200,200,201,202,202,203,204,205,205,206,207,207,208,209,209,210,211,212,212,213,214,214,215,216,216,217,218,218,219,220,220,221,222,222,223,224,224,225,226,226,227,228,228,229,230,230,231,232,232,233,234,234,235,235,236,237,237,238,239,239,240,241,241,242,242,243,244,244,245,246,246,247,247,248,249,249,250,251,251,252,252,253,254,254,255,255),
(0,9,13,17,20,23,26,28,30,33,35,37,39,41,43,45,47,48,50,52,53,55,57,58,60,61,63,64,66,67,68,70,71,72,74,75,76,78,79,80,82,83,84,85,87,88,89,90,91,92,94,95,96,97,98,99,100,101,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,165,165,166,167,168,169,169,170,171,172,173,173,174,175,176,176,177,178,179,180,180,181,182,183,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,197,198,199,200,200,201,202,203,203,204,205,205,206,207,207,208,209,210,210,211,212,212,213,214,214,215,216,217,217,218,219,219,220,221,221,222,223,223,224,225,225,226,227,227,228,229,229,230,231,231,232,233,233,234,235,235,236,237,237,238,238,239,240,240,241,242,242,243,244,244,245,245,246,247,247,248,249,249,250,251,251,252,252,253,254,254,255,255),
(0,8,13,16,19,22,25,27,30,32,34,36,38,40,42,44,45,47,49,51,52,54,55,57,58,60,61,63,64,66,67,69,70,71,73,74,75,77,78,79,80,82,83,84,85,86,88,89,90,91,92,93,95,96,97,98,99,100,101,102,103,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,130,131,132,133,134,135,136,137,138,139,140,141,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,154,155,156,157,158,159,159,160,161,162,163,164,164,165,166,167,168,168,169,170,171,172,172,173,174,175,176,176,177,178,179,180,180,181,182,183,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,198,198,199,200,200,201,202,203,203,204,205,205,206,207,208,208,209,210,210,211,212,213,213,214,215,215,216,217,217,218,219,219,220,221,222,222,223,224,224,225,226,226,227,228,228,229,230,230,231,232,232,233,234,234,235,236,236,237,238,238,239,240,240,241,241,242,243,243,244,245,245,246,247,247,248,249,249,250,250,251,252,252,253,254,254,255,255),
(0,8,12,16,19,21,24,26,29,31,33,35,37,39,41,43,44,46,48,50,51,53,54,56,57,59,60,62,63,65,66,67,69,70,71,73,74,75,77,78,79,80,82,83,84,85,86,88,89,90,91,92,93,95,96,97,98,99,100,101,102,103,104,105,106,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,126,127,128,129,130,131,132,133,134,135,136,137,138,139,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,158,159,160,161,162,163,163,164,165,166,167,168,168,169,170,171,172,172,173,174,175,176,176,177,178,179,179,180,181,182,183,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,198,198,199,200,201,201,202,203,203,204,205,206,206,207,208,208,209,210,211,211,212,213,213,214,215,216,216,217,218,218,219,220,220,221,222,222,223,224,225,225,226,227,227,228,229,229,230,231,231,232,233,233,234,235,235,236,237,237,238,239,239,240,241,241,242,243,243,244,245,245,246,247,247,248,248,249,250,250,251,252,252,253,254,254,255,255),
(0,8,12,15,18,21,23,26,28,30,32,34,36,38,40,42,43,45,47,48,50,52,53,55,56,58,59,61,62,63,65,66,68,69,70,72,73,74,75,77,78,79,80,82,83,84,85,86,88,89,90,91,92,93,94,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,116,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,136,137,138,139,140,141,142,143,144,145,145,146,147,148,149,150,151,152,152,153,154,155,156,157,157,158,159,160,161,162,162,163,164,165,166,167,167,168,169,170,171,171,172,173,174,175,175,176,177,178,179,179,180,181,182,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,198,198,199,200,201,201,202,203,204,204,205,206,206,207,208,209,209,210,211,212,212,213,214,214,215,216,216,217,218,219,219,220,221,221,222,223,223,224,225,226,226,227,228,228,229,230,230,231,232,232,233,234,234,235,236,236,237,238,238,239,240,240,241,242,242,243,244,244,245,246,246,247,248,248,249,250,250,251,252,252,253,254,254,255,255),
(0,7,11,15,17,20,23,25,27,29,31,33,35,37,39,41,42,44,46,47,49,51,52,54,55,57,58,59,61,62,64,65,66,68,69,70,72,73,74,75,77,78,79,80,82,83,84,85,86,87,89,90,91,92,93,94,95,96,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,150,151,152,153,154,155,156,156,157,158,159,160,161,161,162,163,164,165,166,166,167,168,169,170,171,171,172,173,174,175,175,176,177,178,179,179,180,181,182,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,195,196,197,198,198,199,200,201,201,202,203,204,204,205,206,207,207,208,209,210,210,211,212,212,213,214,215,215,216,217,217,218,219,220,220,221,222,222,223,224,224,225,226,227,227,228,229,229,230,231,231,232,233,233,234,235,236,236,237,238,238,239,240,240,241,242,242,243,244,244,245,246,246,247,248,248,249,250,250,251,252,252,253,254,254,255,255),
(0,7,11,14,17,19,22,24,26,28,30,32,34,36,38,40,41,43,45,46,48,49,51,52,54,55,57,58,60,61,62,64,65,66,68,69,70,72,73,74,75,77,78,79,80,81,83,84,85,86,87,88,90,91,92,93,94,95,96,97,98,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,130,131,132,133,134,135,136,137,138,139,140,141,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,155,155,156,157,158,159,160,160,161,162,163,164,165,165,166,167,168,169,170,170,171,172,173,174,174,175,176,177,178,178,179,180,181,182,182,183,184,185,186,186,187,188,189,189,190,191,192,192,193,194,195,196,196,197,198,199,199,200,201,202,202,203,204,205,205,206,207,207,208,209,210,210,211,212,213,213,214,215,215,216,217,218,218,219,220,221,221,222,223,223,224,225,225,226,227,228,228,229,230,230,231,232,232,233,234,235,235,236,237,237,238,239,239,240,241,241,242,243,243,244,245,245,246,247,248,248,249,250,250,251,252,252,253,254,254,255,255),
(0,7,10,13,16,19,21,23,26,28,30,32,33,35,37,39,40,42,44,45,47,48,50,51,53,54,56,57,58,60,61,63,64,65,67,68,69,70,72,73,74,75,77,78,79,80,81,83,84,85,86,87,88,89,91,92,93,94,95,96,97,98,99,100,101,102,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,125,126,127,128,129,130,131,132,133,134,135,136,137,138,138,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,153,154,155,156,157,158,159,159,160,161,162,163,164,164,165,166,167,168,169,169,170,171,172,173,174,174,175,176,177,178,178,179,180,181,182,182,183,184,185,186,186,187,188,189,189,190,191,192,193,193,194,195,196,196,197,198,199,199,200,201,202,202,203,204,205,205,206,207,208,208,209,210,211,211,212,213,214,214,215,216,216,217,218,219,219,220,221,222,222,223,224,224,225,226,227,227,228,229,229,230,231,231,232,233,234,234,235,236,236,237,238,238,239,240,241,241,242,243,243,244,245,245,246,247,247,248,249,249,250,251,251,252,253,253,254,255,255),
(0,6,10,13,16,18,20,23,25,27,29,31,32,34,36,38,39,41,43,44,46,47,49,50,52,53,55,56,57,59,60,61,63,64,65,67,68,69,70,72,73,74,75,77,78,79,80,81,82,84,85,86,87,88,89,90,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,113,114,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,135,136,137,138,139,140,141,142,143,144,145,145,146,147,148,149,150,151,152,152,153,154,155,156,157,158,158,159,160,161,162,163,163,164,165,166,167,168,168,169,170,171,172,173,173,174,175,176,177,177,178,179,180,181,182,182,183,184,185,185,186,187,188,189,189,190,191,192,193,193,194,195,196,196,197,198,199,199,200,201,202,203,203,204,205,206,206,207,208,209,209,210,211,212,212,213,214,214,215,216,217,217,218,219,220,220,221,222,223,223,224,225,225,226,227,228,228,229,230,230,231,232,233,233,234,235,235,236,237,238,238,239,240,240,241,242,242,243,244,245,245,246,247,247,248,249,249,250,251,251,252,253,253,254,255,255),
(0,6,10,12,15,17,20,22,24,26,28,30,32,33,35,37,38,40,42,43,45,46,48,49,51,52,53,55,56,58,59,60,62,63,64,65,67,68,69,70,72,73,74,75,76,78,79,80,81,82,83,85,86,87,88,89,90,91,92,93,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,131,132,133,134,135,136,137,138,139,140,141,142,142,143,144,145,146,147,148,149,150,150,151,152,153,154,155,156,157,157,158,159,160,161,162,162,163,164,165,166,167,168,168,169,170,171,172,172,173,174,175,176,177,177,178,179,180,181,181,182,183,184,185,185,186,187,188,189,189,190,191,192,193,193,194,195,196,196,197,198,199,200,200,201,202,203,203,204,205,206,206,207,208,209,209,210,211,212,212,213,214,215,215,216,217,218,218,219,220,221,221,222,223,224,224,225,226,226,227,228,229,229,230,231,232,232,233,234,234,235,236,237,237,238,239,239,240,241,242,242,243,244,244,245,246,246,247,248,249,249,250,251,251,252,253,253,254,255,255),
(0,6,9,12,14,17,19,21,23,25,27,29,31,32,34,36,37,39,40,42,44,45,47,48,49,51,52,54,55,56,58,59,60,62,63,64,65,67,68,69,70,72,73,74,75,76,78,79,80,81,82,83,84,86,87,88,89,90,91,92,93,94,95,96,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,127,128,129,130,131,132,133,134,135,136,137,138,139,139,140,141,142,143,144,145,146,147,148,148,149,150,151,152,153,154,155,155,156,157,158,159,160,161,161,162,163,164,165,166,167,167,168,169,170,171,172,172,173,174,175,176,176,177,178,179,180,181,181,182,183,184,185,185,186,187,188,189,189,190,191,192,193,193,194,195,196,197,197,198,199,200,200,201,202,203,204,204,205,206,207,207,208,209,210,210,211,212,213,213,214,215,216,216,217,218,219,219,220,221,222,222,223,224,225,225,226,227,228,228,229,230,231,231,232,233,233,234,235,236,236,237,238,238,239,240,241,241,242,243,243,244,245,246,246,247,248,248,249,250,251,251,252,253,253,254,255,255),
(0,6,9,11,14,16,18,20,22,24,26,28,30,31,33,35,36,38,39,41,42,44,45,47,48,50,51,52,54,55,56,58,59,60,62,63,64,65,67,68,69,70,72,73,74,75,76,77,79,80,81,82,83,84,85,86,88,89,90,91,92,93,94,95,96,97,98,99,100,101,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,136,137,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,153,153,154,155,156,157,158,159,160,160,161,162,163,164,165,166,166,167,168,169,170,171,171,172,173,174,175,176,176,177,178,179,180,181,181,182,183,184,185,185,186,187,188,189,189,190,191,192,193,193,194,195,196,197,197,198,199,200,201,201,202,203,204,204,205,206,207,207,208,209,210,211,211,212,213,214,214,215,216,217,217,218,219,220,220,221,222,223,223,224,225,226,226,227,228,229,229,230,231,232,232,233,234,235,235,236,237,238,238,239,240,240,241,242,243,243,244,245,245,246,247,248,248,249,250,251,251,252,253,253,254,255,255),
(0,5,8,11,13,16,18,20,22,24,25,27,29,31,32,34,35,37,38,40,41,43,44,46,47,49,50,51,53,54,55,57,58,59,60,62,63,64,65,67,68,69,70,71,73,74,75,76,77,78,80,81,82,83,84,85,86,87,88,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,132,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,151,151,152,153,154,155,156,157,158,158,159,160,161,162,163,164,164,165,166,167,168,169,170,170,171,172,173,174,175,175,176,177,178,179,180,180,181,182,183,184,185,185,186,187,188,189,189,190,191,192,193,193,194,195,196,197,197,198,199,200,201,201,202,203,204,205,205,206,207,208,208,209,210,211,212,212,213,214,215,215,216,217,218,218,219,220,221,222,222,223,224,225,225,226,227,228,228,229,230,231,231,232,233,234,234,235,236,237,237,238,239,239,240,241,242,242,243,244,245,245,246,247,248,248,249,250,250,251,252,253,253,254,255,255),
(0,5,8,10,13,15,17,19,21,23,25,26,28,30,31,33,34,36,37,39,40,42,43,45,46,47,49,50,51,53,54,55,57,58,59,60,62,63,64,65,67,68,69,70,71,72,74,75,76,77,78,79,80,82,83,84,85,86,87,88,89,90,91,92,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,127,128,129,130,131,132,133,134,135,136,137,138,139,140,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,156,157,157,158,159,160,161,162,163,163,164,165,166,167,168,169,169,170,171,172,173,174,175,175,176,177,178,179,180,180,181,182,183,184,184,185,186,187,188,189,189,190,191,192,193,193,194,195,196,197,197,198,199,200,201,201,202,203,204,205,205,206,207,208,209,209,210,211,212,213,213,214,215,216,216,217,218,219,220,220,221,222,223,223,224,225,226,226,227,228,229,229,230,231,232,232,233,234,235,236,236,237,238,239,239,240,241,241,242,243,244,244,245,246,247,247,248,249,250,250,251,252,253,253,254,255,255),
(0,5,8,10,12,14,16,18,20,22,24,25,27,29,30,32,33,35,36,38,39,41,42,44,45,46,48,49,50,52,53,54,55,57,58,59,60,62,63,64,65,66,68,69,70,71,72,73,75,76,77,78,79,80,81,82,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,136,137,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,161,162,162,163,164,165,166,167,168,168,169,170,171,172,173,174,174,175,176,177,178,179,179,180,181,182,183,184,184,185,186,187,188,189,189,190,191,192,193,194,194,195,196,197,198,198,199,200,201,202,202,203,204,205,206,206,207,208,209,210,210,211,212,213,214,214,215,216,217,217,218,219,220,221,221,222,223,224,224,225,226,227,228,228,229,230,231,231,232,233,234,234,235,236,237,238,238,239,240,241,241,242,243,244,244,245,246,247,247,248,249,250,250,251,252,253,253,254,255,255),
(0,4,7,10,12,14,16,18,19,21,23,25,26,28,29,31,32,34,35,37,38,40,41,42,44,45,46,48,49,50,52,53,54,55,57,58,59,60,62,63,64,65,66,68,69,70,71,72,73,74,76,77,78,79,80,81,82,83,84,85,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,131,132,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,151,152,152,153,154,155,156,157,158,159,160,160,161,162,163,164,165,166,167,167,168,169,170,171,172,173,173,174,175,176,177,178,179,179,180,181,182,183,184,184,185,186,187,188,189,189,190,191,192,193,194,194,195,196,197,198,198,199,200,201,202,203,203,204,205,206,207,207,208,209,210,211,211,212,213,214,215,215,216,217,218,219,219,220,221,222,222,223,224,225,226,226,227,228,229,230,230,231,232,233,233,234,235,236,236,237,238,239,240,240,241,242,243,243,244,245,246,246,247,248,249,249,250,251,252,252,253,254,255,255),
(0,4,7,9,11,13,15,17,19,20,22,24,25,27,28,30,31,33,34,36,37,39,40,41,43,44,45,47,48,49,50,52,53,54,55,57,58,59,60,61,63,64,65,66,67,69,70,71,72,73,74,75,76,78,79,80,81,82,83,84,85,86,87,88,89,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,140,141,142,143,144,145,146,147,148,149,150,150,151,152,153,154,155,156,157,158,158,159,160,161,162,163,164,165,165,166,167,168,169,170,171,172,172,173,174,175,176,177,178,178,179,180,181,182,183,184,184,185,186,187,188,189,189,190,191,192,193,194,194,195,196,197,198,199,199,200,201,202,203,203,204,205,206,207,208,208,209,210,211,212,212,213,214,215,216,216,217,218,219,220,220,221,222,223,224,224,225,226,227,228,228,229,230,231,232,232,233,234,235,235,236,237,238,239,239,240,241,242,242,243,244,245,246,246,247,248,249,249,250,251,252,252,253,254,255,255),
(0,4,7,9,11,13,15,16,18,20,21,23,24,26,28,29,30,32,33,35,36,37,39,40,42,43,44,45,47,48,49,50,52,53,54,55,57,58,59,60,61,63,64,65,66,67,68,69,71,72,73,74,75,76,77,78,79,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,101,102,103,104,105,106,107,108,109,110,111,112,113,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,135,136,137,138,139,140,141,142,143,144,145,146,147,147,148,149,150,151,152,153,154,155,156,156,157,158,159,160,161,162,163,164,164,165,166,167,168,169,170,171,171,172,173,174,175,176,177,177,178,179,180,181,182,183,183,184,185,186,187,188,189,189,190,191,192,193,194,194,195,196,197,198,199,199,200,201,202,203,204,204,205,206,207,208,209,209,210,211,212,213,213,214,215,216,217,218,218,219,220,221,222,222,223,224,225,226,226,227,228,229,230,230,231,232,233,234,234,235,236,237,238,238,239,240,241,241,242,243,244,245,245,246,247,248,249,249,250,251,252,252,253,254,255,255),
(0,4,6,8,10,12,14,16,17,19,21,22,24,25,27,28,30,31,32,34,35,36,38,39,40,42,43,44,46,47,48,49,51,52,53,54,55,57,58,59,60,61,62,64,65,66,67,68,69,70,71,73,74,75,76,77,78,79,80,81,82,83,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,143,144,145,146,147,148,149,150,151,152,153,153,154,155,156,157,158,159,160,161,162,162,163,164,165,166,167,168,169,170,170,171,172,173,174,175,176,177,177,178,179,180,181,182,183,183,184,185,186,187,188,189,189,190,191,192,193,194,195,195,196,197,198,199,200,200,201,202,203,204,205,205,206,207,208,209,210,210,211,212,213,214,215,215,216,217,218,219,219,220,221,222,223,224,224,225,226,227,228,228,229,230,231,232,232,233,234,235,236,236,237,238,239,240,240,241,242,243,244,244,245,246,247,248,248,249,250,251,252,252,253,254,255,255),
(0,4,6,8,10,12,13,15,17,18,20,21,23,24,26,27,29,30,31,33,34,35,37,38,39,41,42,43,44,46,47,48,49,50,52,53,54,55,56,58,59,60,61,62,63,65,66,67,68,69,70,71,72,73,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,138,139,140,141,142,143,144,145,146,147,148,149,150,150,151,152,153,154,155,156,157,158,159,160,160,161,162,163,164,165,166,167,168,168,169,170,171,172,173,174,175,176,176,177,178,179,180,181,182,182,183,184,185,186,187,188,189,189,190,191,192,193,194,195,195,196,197,198,199,200,201,201,202,203,204,205,206,206,207,208,209,210,211,211,212,213,214,215,216,216,217,218,219,220,221,221,222,223,224,225,226,226,227,228,229,230,230,231,232,233,234,235,235,236,237,238,239,239,240,241,242,243,243,244,245,246,247,247,248,249,250,251,252,252,253,254,255,255),
(0,3,6,8,9,11,13,14,16,18,19,21,22,23,25,26,28,29,30,32,33,34,36,37,38,39,41,42,43,44,46,47,48,49,50,52,53,54,55,56,57,59,60,61,62,63,64,65,67,68,69,70,71,72,73,74,75,76,77,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,153,154,155,156,157,157,158,159,160,161,162,163,164,165,166,166,167,168,169,170,171,172,173,174,175,175,176,177,178,179,180,181,182,182,183,184,185,186,187,188,189,189,190,191,192,193,194,195,195,196,197,198,199,200,201,201,202,203,204,205,206,207,207,208,209,210,211,212,213,213,214,215,216,217,218,218,219,220,221,222,223,223,224,225,226,227,228,228,229,230,231,232,233,233,234,235,236,237,238,238,239,240,241,242,242,243,244,245,246,247,247,248,249,250,251,251,252,253,254,255,255),
(0,3,5,7,9,11,12,14,15,17,18,20,21,23,24,25,27,28,29,31,32,33,35,36,37,38,40,41,42,43,44,46,47,48,49,50,52,53,54,55,56,57,58,60,61,62,63,64,65,66,67,68,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,142,143,144,145,146,147,148,149,150,151,152,153,154,154,155,156,157,158,159,160,161,162,163,164,164,165,166,167,168,169,170,171,172,173,173,174,175,176,177,178,179,180,181,181,182,183,184,185,186,187,188,189,189,190,191,192,193,194,195,196,196,197,198,199,200,201,202,202,203,204,205,206,207,208,208,209,210,211,212,213,214,214,215,216,217,218,219,220,220,221,222,223,224,225,226,226,227,228,229,230,231,231,232,233,234,235,236,236,237,238,239,240,241,241,242,243,244,245,246,246,247,248,249,250,251,251,252,253,254,255,255),
(0,3,5,7,8,10,12,13,15,16,18,19,20,22,23,24,26,27,28,30,31,32,33,35,36,37,38,40,41,42,43,44,46,47,48,49,50,51,53,54,55,56,57,58,59,60,62,63,64,65,66,67,68,69,70,71,72,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,150,151,152,153,154,155,156,157,158,159,160,161,162,162,163,164,165,166,167,168,169,170,171,172,172,173,174,175,176,177,178,179,180,181,181,182,183,184,185,186,187,188,189,189,190,191,192,193,194,195,196,196,197,198,199,200,201,202,203,203,204,205,206,207,208,209,210,210,211,212,213,214,215,216,216,217,218,219,220,221,222,223,223,224,225,226,227,228,229,229,230,231,232,233,234,234,235,236,237,238,239,240,240,241,242,243,244,245,245,246,247,248,249,250,250,251,252,253,254,255,255),
(0,3,5,6,8,10,11,13,14,15,17,18,20,21,22,24,25,26,27,29,30,31,32,34,35,36,37,39,40,41,42,43,44,46,47,48,49,50,51,52,54,55,56,57,58,59,60,61,62,63,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,159,160,161,162,163,164,165,166,167,168,169,170,170,171,172,173,174,175,176,177,178,179,180,180,181,182,183,184,185,186,187,188,189,189,190,191,192,193,194,195,196,197,197,198,199,200,201,202,203,204,205,205,206,207,208,209,210,211,212,212,213,214,215,216,217,218,219,219,220,221,222,223,224,225,226,226,227,228,229,230,231,232,232,233,234,235,236,237,238,238,239,240,241,242,243,244,244,245,246,247,248,249,250,250,251,252,253,254,255,255),
(0,3,4,6,8,9,11,12,13,15,16,18,19,20,21,23,24,25,26,28,29,30,31,33,34,35,36,37,39,40,41,42,43,44,45,47,48,49,50,51,52,53,54,56,57,58,59,60,61,62,63,64,65,66,67,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,161,162,163,164,165,166,167,168,168,169,170,171,172,173,174,175,176,177,178,179,179,180,181,182,183,184,185,186,187,188,189,189,190,191,192,193,194,195,196,197,198,198,199,200,201,202,203,204,205,206,206,207,208,209,210,211,212,213,214,214,215,216,217,218,219,220,221,222,222,223,224,225,226,227,228,229,229,230,231,232,233,234,235,236,236,237,238,239,240,241,242,243,243,244,245,246,247,248,249,249,250,251,252,253,254,255,255),
(0,2,4,6,7,9,10,11,13,14,15,17,18,19,21,22,23,24,26,27,28,29,30,32,33,34,35,36,37,39,40,41,42,43,44,45,46,48,49,50,51,52,53,54,55,56,57,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,165,166,167,168,169,170,171,172,173,174,175,176,177,177,178,179,180,181,182,183,184,185,186,187,188,188,189,190,191,192,193,194,195,196,197,198,199,199,200,201,202,203,204,205,206,207,208,208,209,210,211,212,213,214,215,216,217,217,218,219,220,221,222,223,224,225,225,226,227,228,229,230,231,232,233,233,234,235,236,237,238,239,240,241,241,242,243,244,245,246,247,248,248,249,250,251,252,253,254,255,255),
(0,2,4,5,7,8,10,11,12,14,15,16,17,19,20,21,22,23,25,26,27,28,29,31,32,33,34,35,36,37,39,40,41,42,43,44,45,46,47,48,50,51,52,53,54,55,56,57,58,59,60,61,62,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,175,176,177,178,179,180,181,182,183,184,185,186,187,188,188,189,190,191,192,193,194,195,196,197,198,199,200,200,201,202,203,204,205,206,207,208,209,210,211,211,212,213,214,215,216,217,218,219,220,220,221,222,223,224,225,226,227,228,229,230,230,231,232,233,234,235,236,237,238,239,239,240,241,242,243,244,245,246,247,247,248,249,250,251,252,253,254,255,255),
(0,2,4,5,6,8,9,10,12,13,14,15,17,18,19,20,21,23,24,25,26,27,28,29,31,32,33,34,35,36,37,38,40,41,42,43,44,45,46,47,48,49,50,51,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,202,203,204,205,206,207,208,209,210,211,212,213,214,214,215,216,217,218,219,220,221,222,223,224,225,225,226,227,228,229,230,231,232,233,234,235,236,236,237,238,239,240,241,242,243,244,245,246,246,247,248,249,250,251,252,253,254,255,255),
(0,2,3,5,6,7,9,10,11,12,13,15,16,17,18,19,21,22,23,24,25,26,27,28,30,31,32,33,34,35,36,37,38,39,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,218,219,220,221,222,223,224,225,226,227,228,229,230,231,231,232,233,234,235,236,237,238,239,240,241,242,243,244,244,245,246,247,248,249,250,251,252,253,254,255,255),
(0,2,3,5,6,7,8,9,11,12,13,14,15,16,17,19,20,21,22,23,24,25,26,27,28,30,31,32,33,34,35,36,37,38,39,40,41,42,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255,255),
(0,2,3,4,5,7,8,9,10,11,12,13,14,16,17,18,19,20,21,22,23,24,25,26,27,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,213,214,215,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255,255),
(0,2,3,4,5,6,7,8,9,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,185,186,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,224,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255,255),
(0,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255,255),
(0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255),
(0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255),
(0,1,2,3,4,5,6,7,8,8,9,10,11,12,13,14,15,16,17,18,19,20,21,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,192,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,226,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255),
(0,1,2,3,4,4,5,6,7,8,9,10,11,11,12,13,14,15,16,17,18,19,20,21,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255),
(0,1,2,3,3,4,5,6,7,7,8,9,10,11,12,13,13,14,15,16,17,18,19,20,21,21,22,23,24,25,26,27,28,29,30,31,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,227,228,229,230,231,232,233,234,235,236,237,238,239,240,242,243,244,245,246,247,248,249,250,251,252,253,254,255),
(0,1,2,2,3,4,5,5,6,7,8,9,9,10,11,12,13,14,14,15,16,17,18,19,20,20,21,22,23,24,25,26,27,28,28,29,30,31,32,33,34,35,36,37,38,39,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,192,193,194,195,196,197,198,199,200,201,202,203,204,205,207,208,209,210,211,212,213,214,215,216,217,218,220,221,222,223,224,225,226,227,228,229,230,231,233,234,235,236,237,238,239,240,241,242,243,245,246,247,248,249,250,251,252,253,254,255),
(0,1,2,2,3,4,4,5,6,7,7,8,9,10,10,11,12,13,14,14,15,16,17,18,19,19,20,21,22,23,24,25,26,26,27,28,29,30,31,32,33,34,34,35,36,37,38,39,40,41,42,43,44,45,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,163,164,165,166,167,168,169,170,171,172,173,174,175,176,178,179,180,181,182,183,184,185,186,187,188,189,190,192,193,194,195,196,197,198,199,200,201,202,204,205,206,207,208,209,210,211,212,213,214,216,217,218,219,220,221,222,223,224,226,227,228,229,230,231,232,233,234,235,237,238,239,240,241,242,243,244,245,247,248,249,250,251,252,253,254,255),
(0,1,2,2,3,3,4,5,5,6,7,8,8,9,10,11,11,12,13,14,15,15,16,17,18,19,19,20,21,22,23,24,24,25,26,27,28,29,30,30,31,32,33,34,35,36,37,38,38,39,40,41,42,43,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,153,154,155,156,157,158,159,160,161,162,163,164,165,167,168,169,170,171,172,173,174,175,176,177,178,180,181,182,183,184,185,186,187,188,189,191,192,193,194,195,196,197,198,199,200,202,203,204,205,206,207,208,209,210,212,213,214,215,216,217,218,219,220,222,223,224,225,226,227,228,229,231,232,233,234,235,236,237,238,240,241,242,243,244,245,246,248,249,250,251,252,253,254,255),
(0,1,1,2,3,3,4,4,5,6,6,7,8,9,9,10,11,11,12,13,14,14,15,16,17,18,18,19,20,21,22,23,23,24,25,26,27,28,28,29,30,31,32,33,34,34,35,36,37,38,39,40,41,42,42,43,44,45,46,47,48,49,50,51,52,53,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,145,146,147,148,149,150,151,152,153,154,155,156,157,159,160,161,162,163,164,165,166,167,168,169,171,172,173,174,175,176,177,178,179,181,182,183,184,185,186,187,188,189,191,192,193,194,195,196,197,198,199,201,202,203,204,205,206,207,208,210,211,212,213,214,215,216,218,219,220,221,222,223,224,226,227,228,229,230,231,232,234,235,236,237,238,239,240,242,243,244,245,246,247,249,250,251,252,253,254,255),
(0,1,1,2,2,3,3,4,5,5,6,7,7,8,9,9,10,11,11,12,13,14,14,15,16,17,18,18,19,20,21,21,22,23,24,25,26,26,27,28,29,30,31,31,32,33,34,35,36,37,37,38,39,40,41,42,43,44,45,45,46,47,48,49,50,51,52,53,54,55,56,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,139,140,141,142,143,144,145,146,147,148,149,150,152,153,154,155,156,157,158,159,160,161,163,164,165,166,167,168,169,170,171,173,174,175,176,177,178,179,180,182,183,184,185,186,187,188,189,191,192,193,194,195,196,197,198,200,201,202,203,204,205,206,208,209,210,211,212,213,215,216,217,218,219,220,221,223,224,225,226,227,228,230,231,232,233,234,235,237,238,239,240,241,243,244,245,246,247,248,250,251,252,253,254,255),
(0,1,1,2,2,3,3,4,4,5,6,6,7,7,8,9,9,10,11,12,12,13,14,14,15,16,17,17,18,19,20,20,21,22,23,24,24,25,26,27,28,28,29,30,31,32,33,33,34,35,36,37,38,39,39,40,41,42,43,44,45,46,47,47,48,49,50,51,52,53,54,55,56,57,58,59,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,133,134,135,136,137,138,139,140,141,142,143,144,146,147,148,149,150,151,152,153,154,156,157,158,159,160,161,162,163,164,166,167,168,169,170,171,172,173,175,176,177,178,179,180,181,183,184,185,186,187,188,189,191,192,193,194,195,196,197,199,200,201,202,203,204,206,207,208,209,210,211,213,214,215,216,217,218,220,221,222,223,224,226,227,228,229,230,232,233,234,235,236,237,239,240,241,242,243,245,246,247,248,249,251,252,253,254,255),
(0,1,1,2,2,2,3,4,4,5,5,6,6,7,8,8,9,10,10,11,12,12,13,14,14,15,16,16,17,18,19,19,20,21,22,22,23,24,25,26,26,27,28,29,30,30,31,32,33,34,35,35,36,37,38,39,40,41,41,42,43,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,59,60,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,129,130,131,132,133,134,135,136,137,138,139,141,142,143,144,145,146,147,148,149,151,152,153,154,155,156,157,158,160,161,162,163,164,165,166,168,169,170,171,172,173,174,176,177,178,179,180,181,182,184,185,186,187,188,189,191,192,193,194,195,196,198,199,200,201,202,204,205,206,207,208,209,211,212,213,214,215,217,218,219,220,221,223,224,225,226,227,229,230,231,232,233,235,236,237,238,240,241,242,243,244,246,247,248,249,251,252,253,254,255),
(0,1,1,1,2,2,3,3,4,4,5,5,6,6,7,8,8,9,10,10,11,11,12,13,13,14,15,16,16,17,18,18,19,20,21,21,22,23,24,24,25,26,27,28,28,29,30,31,32,32,33,34,35,36,37,37,38,39,40,41,42,43,43,44,45,46,47,48,49,50,50,51,52,53,54,55,56,57,58,59,60,61,62,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,125,126,127,128,129,130,131,132,133,134,136,137,138,139,140,141,142,143,144,146,147,148,149,150,151,152,153,155,156,157,158,159,160,161,163,164,165,166,167,168,169,171,172,173,174,175,176,178,179,180,181,182,184,185,186,187,188,189,191,192,193,194,195,197,198,199,200,201,203,204,205,206,207,209,210,211,212,213,215,216,217,218,219,221,222,223,224,226,227,228,229,231,232,233,234,235,237,238,239,240,242,243,244,245,247,248,249,250,252,253,254,255),
(0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,7,8,8,9,10,10,11,11,12,13,13,14,15,15,16,17,17,18,19,20,20,21,22,22,23,24,25,26,26,27,28,29,29,30,31,32,33,33,34,35,36,37,38,38,39,40,41,42,43,44,44,45,46,47,48,49,50,51,51,52,53,54,55,56,57,58,59,60,61,62,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,107,108,109,110,111,112,113,114,115,116,117,118,119,120,122,123,124,125,126,127,128,129,130,131,133,134,135,136,137,138,139,140,142,143,144,145,146,147,148,150,151,152,153,154,155,156,158,159,160,161,162,163,165,166,167,168,169,170,172,173,174,175,176,177,179,180,181,182,183,185,186,187,188,189,191,192,193,194,195,197,198,199,200,202,203,204,205,206,208,209,210,211,213,214,215,216,218,219,220,221,223,224,225,226,228,229,230,231,233,234,235,236,238,239,240,241,243,244,245,247,248,249,250,252,253,254,255),
(0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,7,8,8,9,9,10,11,11,12,13,13,14,14,15,16,16,17,18,19,19,20,21,21,22,23,24,24,25,26,27,27,28,29,30,30,31,32,33,34,34,35,36,37,38,39,39,40,41,42,43,44,44,45,46,47,48,49,50,51,51,52,53,54,55,56,57,58,59,60,61,62,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,105,106,107,108,109,110,111,112,113,114,115,116,117,119,120,121,122,123,124,125,126,127,128,130,131,132,133,134,135,136,137,139,140,141,142,143,144,145,147,148,149,150,151,152,154,155,156,157,158,159,161,162,163,164,165,167,168,169,170,171,172,174,175,176,177,178,180,181,182,183,185,186,187,188,189,191,192,193,194,196,197,198,199,201,202,203,204,205,207,208,209,210,212,213,214,216,217,218,219,221,222,223,224,226,227,228,230,231,232,233,235,236,237,239,240,241,242,244,245,246,248,249,250,252,253,254,255),
(0,1,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,7,8,8,9,9,10,11,11,12,12,13,14,14,15,16,16,17,17,18,19,20,20,21,22,22,23,24,25,25,26,27,28,28,29,30,31,31,32,33,34,35,35,36,37,38,39,39,40,41,42,43,44,44,45,46,47,48,49,50,51,51,52,53,54,55,56,57,58,59,60,61,62,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,103,104,105,106,107,108,109,110,111,112,113,114,115,117,118,119,120,121,122,123,124,125,127,128,129,130,131,132,133,134,136,137,138,139,140,141,143,144,145,146,147,148,150,151,152,153,154,155,157,158,159,160,161,163,164,165,166,167,169,170,171,172,173,175,176,177,178,180,181,182,183,184,186,187,188,189,191,192,193,194,196,197,198,199,201,202,203,204,206,207,208,210,211,212,213,215,216,217,219,220,221,222,224,225,226,228,229,230,232,233,234,236,237,238,239,241,242,243,245,246,247,249,250,251,253,254,255),
(0,1,1,1,1,2,2,2,3,3,3,4,4,5,5,6,6,7,7,8,8,9,9,10,10,11,12,12,13,13,14,15,15,16,16,17,18,18,19,20,20,21,22,23,23,24,25,25,26,27,28,28,29,30,31,31,32,33,34,35,35,36,37,38,39,39,40,41,42,43,44,44,45,46,47,48,49,50,51,51,52,53,54,55,56,57,58,59,60,61,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,102,103,104,105,106,107,108,109,110,111,112,113,115,116,117,118,119,120,121,122,123,125,126,127,128,129,130,131,133,134,135,136,137,138,140,141,142,143,144,145,147,148,149,150,151,152,154,155,156,157,158,160,161,162,163,165,166,167,168,169,171,172,173,174,176,177,178,179,181,182,183,184,186,187,188,189,191,192,193,194,196,197,198,200,201,202,203,205,206,207,209,210,211,213,214,215,217,218,219,220,222,223,224,226,227,228,230,231,232,234,235,236,238,239,241,242,243,245,246,247,249,250,251,253,254,255),
(0,1,1,1,1,2,2,2,2,3,3,4,4,4,5,5,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,14,14,15,16,16,17,17,18,19,19,20,21,21,22,23,23,24,25,26,26,27,28,29,29,30,31,32,32,33,34,35,35,36,37,38,39,39,40,41,42,43,44,44,45,46,47,48,49,50,50,51,52,53,54,55,56,57,58,59,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,102,103,104,105,106,107,108,109,110,111,112,114,115,116,117,118,119,120,121,123,124,125,126,127,128,129,131,132,133,134,135,136,138,139,140,141,142,144,145,146,147,148,149,151,152,153,154,156,157,158,159,160,162,163,164,165,167,168,169,170,172,173,174,175,177,178,179,180,182,183,184,186,187,188,189,191,192,193,195,196,197,198,200,201,202,204,205,206,208,209,210,212,213,214,216,217,218,220,221,222,224,225,226,228,229,231,232,233,235,236,237,239,240,242,243,244,246,247,248,250,251,253,254,255),
(0,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,15,15,16,16,17,18,18,19,20,20,21,22,22,23,24,24,25,26,26,27,28,29,29,30,31,32,32,33,34,35,35,36,37,38,39,39,40,41,42,43,44,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,102,103,104,105,106,107,108,109,110,111,113,114,115,116,117,118,119,121,122,123,124,125,126,127,129,130,131,132,133,134,136,137,138,139,140,142,143,144,145,146,148,149,150,151,153,154,155,156,157,159,160,161,162,164,165,166,167,169,170,171,173,174,175,176,178,179,180,182,183,184,185,187,188,189,191,192,193,195,196,197,199,200,201,203,204,205,207,208,209,211,212,213,215,216,218,219,220,222,223,224,226,227,229,230,231,233,234,236,237,238,240,241,243,244,245,247,248,250,251,253,254,255),
(0,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,12,12,13,14,14,15,15,16,17,17,18,18,19,20,20,21,22,22,23,24,24,25,26,26,27,28,29,29,30,31,32,32,33,34,35,35,36,37,38,38,39,40,41,42,43,43,44,45,46,47,48,48,49,50,51,52,53,54,55,56,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,71,72,73,74,75,76,77,78,79,80,81,82,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,102,103,104,105,106,107,108,109,110,112,113,114,115,116,117,118,120,121,122,123,124,125,127,128,129,130,131,132,134,135,136,137,138,140,141,142,143,145,146,147,148,149,151,152,153,154,156,157,158,159,161,162,163,165,166,167,168,170,171,172,174,175,176,177,179,180,181,183,184,185,187,188,189,191,192,193,195,196,197,199,200,202,203,204,206,207,208,210,211,213,214,215,217,218,220,221,222,224,225,227,228,229,231,232,234,235,237,238,239,241,242,244,245,247,248,250,251,253,254,255),
(0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15,16,16,17,17,18,19,19,20,20,21,22,22,23,24,24,25,26,26,27,28,29,29,30,31,31,32,33,34,34,35,36,37,38,38,39,40,41,42,42,43,44,45,46,47,47,48,49,50,51,52,53,54,54,55,56,57,58,59,60,61,62,63,64,65,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,88,89,90,91,92,93,94,95,96,97,98,99,100,102,103,104,105,106,107,108,109,110,112,113,114,115,116,117,119,120,121,122,123,124,126,127,128,129,130,132,133,134,135,136,138,139,140,141,143,144,145,146,148,149,150,151,153,154,155,156,158,159,160,162,163,164,165,167,168,169,171,172,173,175,176,177,179,180,181,183,184,185,187,188,189,191,192,194,195,196,198,199,200,202,203,205,206,207,209,210,212,213,214,216,217,219,220,222,223,225,226,227,229,230,232,233,235,236,238,239,241,242,244,245,247,248,249,251,252,254,255),
(0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,8,9,9,10,10,11,11,12,12,13,13,14,15,15,16,16,17,17,18,19,19,20,20,21,22,22,23,24,24,25,26,26,27,28,28,29,30,31,31,32,33,34,34,35,36,37,37,38,39,40,41,41,42,43,44,45,46,46,47,48,49,50,51,52,52,53,54,55,56,57,58,59,60,61,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,91,92,93,94,95,96,97,98,99,100,101,103,104,105,106,107,108,109,111,112,113,114,115,116,117,119,120,121,122,123,125,126,127,128,129,131,132,133,134,136,137,138,139,141,142,143,144,146,147,148,149,151,152,153,155,156,157,158,160,161,162,164,165,166,168,169,170,172,173,174,176,177,178,180,181,183,184,185,187,188,189,191,192,194,195,196,198,199,201,202,203,205,206,208,209,211,212,214,215,216,218,219,221,222,224,225,227,228,230,231,233,234,236,237,239,240,242,243,245,246,248,249,251,252,254,255),
(0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,10,11,11,12,12,13,14,14,15,15,16,16,17,17,18,19,19,20,20,21,22,22,23,24,24,25,26,26,27,28,28,29,30,30,31,32,33,33,34,35,36,36,37,38,39,40,40,41,42,43,44,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,93,94,95,96,97,98,99,100,101,103,104,105,106,107,108,109,111,112,113,114,115,116,118,119,120,121,122,124,125,126,127,128,130,131,132,133,135,136,137,138,140,141,142,144,145,146,147,149,150,151,153,154,155,157,158,159,161,162,163,165,166,167,169,170,171,173,174,175,177,178,180,181,182,184,185,187,188,189,191,192,194,195,197,198,199,201,202,204,205,207,208,210,211,213,214,216,217,219,220,222,223,225,226,228,229,231,232,234,235,237,238,240,241,243,245,246,248,249,251,252,254,255),
(0,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,19,19,20,20,21,22,22,23,24,24,25,25,26,27,27,28,29,30,30,31,32,32,33,34,35,35,36,37,38,39,39,40,41,42,42,43,44,45,46,47,47,48,49,50,51,52,53,54,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,68,69,70,71,72,73,74,75,76,77,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,95,96,97,98,99,100,101,102,104,105,106,107,108,109,111,112,113,114,115,116,118,119,120,121,123,124,125,126,127,129,130,131,132,134,135,136,138,139,140,141,143,144,145,147,148,149,151,152,153,155,156,157,159,160,161,163,164,165,167,168,170,171,172,174,175,177,178,179,181,182,184,185,187,188,189,191,192,194,195,197,198,200,201,203,204,206,207,209,210,212,213,215,216,218,219,221,222,224,225,227,228,230,232,233,235,236,238,239,241,243,244,246,247,249,251,252,254,255),
(0,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,19,19,20,20,21,21,22,23,23,24,25,25,26,27,27,28,29,29,30,31,31,32,33,34,34,35,36,37,37,38,39,40,41,41,42,43,44,45,45,46,47,48,49,50,51,51,52,53,54,55,56,57,58,59,60,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,85,86,87,88,89,90,91,92,93,94,95,97,98,99,100,101,102,103,105,106,107,108,109,111,112,113,114,115,117,118,119,120,121,123,124,125,126,128,129,130,131,133,134,135,137,138,139,141,142,143,145,146,147,149,150,151,153,154,155,157,158,159,161,162,164,165,166,168,169,171,172,173,175,176,178,179,181,182,184,185,186,188,189,191,192,194,195,197,198,200,201,203,204,206,207,209,211,212,214,215,217,218,220,221,223,225,226,228,229,231,233,234,236,237,239,241,242,244,246,247,249,251,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,20,20,21,21,22,23,23,24,24,25,26,26,27,28,28,29,30,30,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,43,43,44,45,46,47,48,48,49,50,51,52,53,54,55,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,89,90,91,92,93,94,95,96,98,99,100,101,102,103,105,106,107,108,109,110,112,113,114,115,117,118,119,120,122,123,124,125,127,128,129,130,132,133,134,136,137,138,140,141,142,144,145,146,148,149,150,152,153,155,156,157,159,160,162,163,164,166,167,169,170,172,173,175,176,177,179,180,182,183,185,186,188,189,191,192,194,195,197,199,200,202,203,205,206,208,209,211,213,214,216,217,219,221,222,224,225,227,229,230,232,234,235,237,239,240,242,244,245,247,249,250,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,21,21,22,22,23,24,24,25,25,26,27,27,28,29,29,30,31,32,32,33,34,34,35,36,37,37,38,39,40,41,41,42,43,44,45,45,46,47,48,49,50,51,51,52,53,54,55,56,57,58,59,60,61,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,80,81,82,83,84,85,86,87,88,89,90,92,93,94,95,96,97,98,100,101,102,103,104,106,107,108,109,110,112,113,114,115,117,118,119,120,122,123,124,126,127,128,129,131,132,133,135,136,137,139,140,141,143,144,146,147,148,150,151,153,154,155,157,158,160,161,162,164,165,167,168,170,171,173,174,176,177,179,180,182,183,185,186,188,189,191,193,194,196,197,199,200,202,204,205,207,208,210,212,213,215,216,218,220,221,223,225,226,228,230,231,233,235,236,238,240,242,243,245,247,249,250,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,5,6,6,6,6,7,7,8,8,8,9,9,9,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,17,18,18,19,19,20,20,21,21,22,23,23,24,25,25,26,26,27,28,28,29,30,30,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,42,43,44,45,46,47,47,48,49,50,51,52,53,54,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,85,86,87,88,89,90,91,92,94,95,96,97,98,99,101,102,103,104,105,107,108,109,110,112,113,114,115,117,118,119,120,122,123,124,126,127,128,130,131,132,134,135,136,138,139,140,142,143,145,146,147,149,150,152,153,155,156,158,159,160,162,163,165,166,168,169,171,172,174,175,177,178,180,182,183,185,186,188,189,191,193,194,196,197,199,201,202,204,206,207,209,210,212,214,215,217,219,221,222,224,226,227,229,231,232,234,236,238,239,241,243,245,247,248,250,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,21,21,22,22,23,24,24,25,25,26,27,27,28,29,29,30,31,31,32,33,34,34,35,36,37,37,38,39,40,40,41,42,43,44,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,59,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,77,78,79,80,81,82,83,84,85,86,88,89,90,91,92,93,94,96,97,98,99,100,102,103,104,105,106,108,109,110,111,113,114,115,117,118,119,120,122,123,124,126,127,128,130,131,133,134,135,137,138,140,141,142,144,145,147,148,150,151,152,154,155,157,158,160,161,163,164,166,167,169,170,172,174,175,177,178,180,181,183,185,186,188,189,191,193,194,196,198,199,201,203,204,206,208,209,211,213,214,216,218,220,221,223,225,227,228,230,232,234,235,237,239,241,243,244,246,248,250,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15,15,16,16,17,18,18,19,19,20,20,21,21,22,23,23,24,24,25,26,26,27,28,28,29,30,30,31,32,32,33,34,35,35,36,37,38,38,39,40,41,41,42,43,44,45,45,46,47,48,49,50,51,52,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,83,84,85,86,87,88,89,91,92,93,94,95,96,98,99,100,101,103,104,105,106,108,109,110,111,113,114,115,117,118,119,121,122,123,125,126,127,129,130,131,133,134,136,137,138,140,141,143,144,146,147,149,150,152,153,155,156,158,159,161,162,164,165,167,168,170,172,173,175,176,178,180,181,183,184,186,188,189,191,193,194,196,198,199,201,203,205,206,208,210,212,213,215,217,219,220,222,224,226,228,229,231,233,235,237,239,240,242,244,246,248,250,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,22,22,23,23,24,25,25,26,26,27,28,28,29,30,30,31,32,33,33,34,35,35,36,37,38,38,39,40,41,42,42,43,44,45,46,47,47,48,49,50,51,52,53,54,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,77,78,79,80,81,82,83,84,85,87,88,89,90,91,92,94,95,96,97,99,100,101,102,104,105,106,107,109,110,111,113,114,115,116,118,119,121,122,123,125,126,127,129,130,132,133,135,136,137,139,140,142,143,145,146,148,149,151,152,154,155,157,158,160,162,163,165,166,168,170,171,173,174,176,178,179,181,183,184,186,188,189,191,193,195,196,198,200,201,203,205,207,209,210,212,214,216,218,219,221,223,225,227,229,231,232,234,236,238,240,242,244,246,248,250,252,254,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,14,15,15,16,16,17,17,18,18,19,19,20,21,21,22,22,23,23,24,25,25,26,27,27,28,29,29,30,31,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,43,43,44,45,46,47,48,48,49,50,51,52,53,54,55,56,57,58,58,59,60,61,62,63,64,65,66,67,68,69,71,72,73,74,75,76,77,78,79,80,81,83,84,85,86,87,88,90,91,92,93,94,96,97,98,99,101,102,103,104,106,107,108,110,111,112,114,115,116,118,119,121,122,123,125,126,128,129,130,132,133,135,136,138,139,141,142,144,145,147,148,150,151,153,155,156,158,159,161,163,164,166,167,169,171,172,174,176,177,179,181,182,184,186,188,189,191,193,195,196,198,200,202,204,205,207,209,211,213,215,217,218,220,222,224,226,228,230,232,234,236,238,240,241,243,245,247,249,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,15,16,16,17,17,18,18,19,20,20,21,21,22,22,23,24,24,25,25,26,27,27,28,29,29,30,31,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,43,43,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,79,80,81,82,83,84,86,87,88,89,90,92,93,94,95,96,98,99,100,102,103,104,105,107,108,109,111,112,114,115,116,118,119,121,122,123,125,126,128,129,131,132,134,135,137,138,140,141,143,144,146,147,149,151,152,154,155,157,159,160,162,164,165,167,169,170,172,174,175,177,179,181,182,184,186,188,189,191,193,195,197,198,200,202,204,206,208,210,212,213,215,217,219,221,223,225,227,229,231,233,235,237,239,241,243,245,247,249,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,22,23,24,24,25,25,26,27,27,28,29,29,30,31,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,43,43,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,75,76,77,78,79,80,81,83,84,85,86,87,89,90,91,92,93,95,96,97,99,100,101,103,104,105,107,108,109,111,112,113,115,116,118,119,120,122,123,125,126,128,129,131,132,134,135,137,138,140,142,143,145,146,148,150,151,153,154,156,158,159,161,163,165,166,168,170,171,173,175,177,179,180,182,184,186,188,189,191,193,195,197,199,201,203,204,206,208,210,212,214,216,218,220,222,224,226,228,230,232,234,236,238,241,243,245,247,249,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,12,13,13,14,14,15,15,16,16,17,17,17,18,19,19,20,20,21,21,22,22,23,23,24,25,25,26,27,27,28,29,29,30,31,31,32,33,33,34,35,36,36,37,38,39,39,40,41,42,43,43,44,45,46,47,48,49,50,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,72,73,74,75,76,77,78,79,81,82,83,84,85,87,88,89,90,92,93,94,95,97,98,99,101,102,103,105,106,108,109,110,112,113,115,116,117,119,120,122,123,125,126,128,129,131,133,134,136,137,139,140,142,144,145,147,149,150,152,154,155,157,159,160,162,164,166,167,169,171,173,175,176,178,180,182,184,186,188,189,191,193,195,197,199,201,203,205,207,209,211,213,215,217,219,221,223,225,227,229,232,234,236,238,240,242,244,247,249,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,8,8,9,9,9,10,10,11,11,11,12,12,12,13,13,14,14,15,15,16,16,16,17,17,18,18,19,19,20,21,21,22,22,23,23,24,25,25,26,26,27,28,28,29,30,30,31,32,32,33,34,35,35,36,37,38,38,39,40,41,42,43,43,44,45,46,47,48,49,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,70,71,72,73,74,75,76,77,79,80,81,82,83,85,86,87,88,90,91,92,94,95,96,98,99,100,102,103,104,106,107,109,110,111,113,114,116,117,119,120,122,123,125,126,128,130,131,133,134,136,138,139,141,142,144,146,148,149,151,153,154,156,158,160,161,163,165,167,169,170,172,174,176,178,180,182,184,186,187,189,191,193,195,197,199,201,203,205,207,210,212,214,216,218,220,222,224,226,229,231,233,235,237,240,242,244,246,249,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,15,16,16,17,17,18,18,19,19,20,20,21,22,22,23,23,24,24,25,26,26,27,28,28,29,30,30,31,32,32,33,34,34,35,36,37,38,38,39,40,41,42,42,43,44,45,46,47,48,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,69,70,71,72,73,74,75,77,78,79,80,81,83,84,85,86,88,89,90,92,93,94,96,97,98,100,101,103,104,105,107,108,110,111,113,114,116,117,119,120,122,123,125,126,128,130,131,133,135,136,138,140,141,143,145,146,148,150,152,153,155,157,159,161,162,164,166,168,170,172,174,176,178,180,181,183,185,187,189,191,193,196,198,200,202,204,206,208,210,212,214,217,219,221,223,225,228,230,232,234,237,239,241,244,246,248,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,22,23,24,24,25,25,26,27,27,28,29,29,30,31,31,32,33,34,34,35,36,37,37,38,39,40,40,41,42,43,44,45,46,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,68,69,70,71,72,73,75,76,77,78,79,81,82,83,84,86,87,88,90,91,92,94,95,96,98,99,101,102,103,105,106,108,109,111,112,114,115,117,118,120,122,123,125,126,128,130,131,133,135,136,138,140,142,143,145,147,149,151,152,154,156,158,160,162,164,165,167,169,171,173,175,177,179,181,183,185,187,189,191,194,196,198,200,202,204,206,209,211,213,215,218,220,222,224,227,229,231,234,236,238,241,243,246,248,251,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,15,16,16,17,17,18,18,19,19,20,20,21,22,22,23,23,24,24,25,26,26,27,28,28,29,30,30,31,32,32,33,34,35,35,36,37,38,39,39,40,41,42,43,44,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,67,68,69,70,71,72,73,75,76,77,78,80,81,82,83,85,86,87,89,90,91,93,94,96,97,98,100,101,103,104,106,107,109,110,112,114,115,117,118,120,122,123,125,126,128,130,132,133,135,137,139,140,142,144,146,148,149,151,153,155,157,159,161,163,165,167,169,171,173,175,177,179,181,183,185,187,189,192,194,196,198,200,203,205,207,209,212,214,216,219,221,223,226,228,231,233,235,238,240,243,245,248,250,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,22,23,24,24,25,25,26,27,27,28,29,29,30,31,31,32,33,34,34,35,36,37,37,38,39,40,41,42,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,68,69,70,71,72,74,75,76,77,79,80,81,82,84,85,87,88,89,91,92,93,95,96,98,99,101,102,104,105,107,108,110,112,113,115,116,118,120,121,123,125,126,128,130,132,133,135,137,139,141,143,144,146,148,150,152,154,156,158,160,162,164,166,168,170,172,174,176,179,181,183,185,187,189,192,194,196,198,201,203,205,208,210,212,215,217,220,222,225,227,230,232,235,237,240,242,245,248,250,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,23,23,24,24,25,26,26,27,27,28,29,30,30,31,32,32,33,34,35,35,36,37,38,39,39,40,41,42,43,44,45,46,46,47,48,49,50,51,52,53,54,55,56,57,59,60,61,62,63,64,65,66,68,69,70,71,72,74,75,76,77,79,80,81,83,84,86,87,88,90,91,93,94,96,97,99,100,102,103,105,106,108,109,111,113,114,116,118,119,121,123,125,126,128,130,132,134,135,137,139,141,143,145,147,149,151,153,155,157,159,161,163,165,167,169,172,174,176,178,180,183,185,187,189,192,194,196,199,201,204,206,208,211,213,216,218,221,223,226,229,231,234,236,239,242,244,247,250,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13,13,14,14,15,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,23,23,24,24,25,26,26,27,28,28,29,30,30,31,32,33,33,34,35,36,36,37,38,39,40,41,42,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,62,63,64,65,66,67,69,70,71,72,74,75,76,78,79,80,82,83,84,86,87,89,90,92,93,95,96,98,99,101,102,104,106,107,109,111,112,114,116,117,119,121,123,125,126,128,130,132,134,136,138,140,142,144,146,148,150,152,154,156,158,160,162,164,167,169,171,173,175,178,180,182,185,187,189,192,194,197,199,202,204,207,209,212,214,217,220,222,225,228,230,233,236,238,241,244,247,250,253,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,6,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,23,23,24,24,25,26,26,27,28,28,29,30,31,31,32,33,33,34,35,36,37,38,38,39,40,41,42,43,44,45,46,46,47,48,49,50,51,52,54,55,56,57,58,59,60,61,62,64,65,66,67,69,70,71,72,74,75,76,78,79,80,82,83,85,86,88,89,91,92,94,95,97,98,100,102,103,105,107,108,110,112,113,115,117,119,121,122,124,126,128,130,132,134,136,138,140,142,144,146,148,150,152,155,157,159,161,163,166,168,170,173,175,177,180,182,184,187,189,192,194,197,200,202,205,207,210,213,215,218,221,224,226,229,232,235,238,241,244,247,249,252,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,23,23,24,24,25,26,26,27,28,28,29,30,31,31,32,33,34,34,35,36,37,38,39,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,59,60,61,62,63,65,66,67,68,70,71,72,74,75,76,78,79,81,82,83,85,86,88,89,91,93,94,96,97,99,101,102,104,106,108,109,111,113,115,117,118,120,122,124,126,128,130,132,134,136,138,140,142,145,147,149,151,153,156,158,160,162,165,167,169,172,174,177,179,182,184,187,189,192,195,197,200,203,205,208,211,214,216,219,222,225,228,231,234,237,240,243,246,249,252,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,22,23,24,24,25,26,26,27,28,28,29,30,31,31,32,33,34,34,35,36,37,38,39,40,40,41,42,43,44,45,46,47,48,49,50,51,52,54,55,56,57,58,59,60,62,63,64,65,67,68,69,71,72,73,75,76,78,79,81,82,84,85,87,88,90,91,93,95,96,98,100,101,103,105,107,109,110,112,114,116,118,120,122,124,126,128,130,132,134,136,138,141,143,145,147,150,152,154,157,159,161,164,166,169,171,174,176,179,181,184,187,189,192,195,198,200,203,206,209,212,215,218,221,224,227,230,233,236,239,242,246,249,252,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17,18,18,19,19,20,21,21,22,22,23,23,24,25,25,26,27,27,28,29,30,30,31,32,33,34,34,35,36,37,38,39,40,41,41,42,43,44,45,46,47,48,50,51,52,53,54,55,56,57,59,60,61,62,64,65,66,68,69,70,72,73,75,76,78,79,81,82,84,85,87,88,90,92,93,95,97,99,100,102,104,106,108,110,112,114,116,118,120,122,124,126,128,130,132,134,137,139,141,143,146,148,150,153,155,158,160,163,165,168,170,173,176,178,181,184,187,189,192,195,198,201,204,207,210,213,216,219,222,225,229,232,235,238,242,245,249,252,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,21,22,23,23,24,24,25,26,27,27,28,29,29,30,31,32,33,33,34,35,36,37,38,39,40,41,41,42,43,44,45,47,48,49,50,51,52,53,54,56,57,58,59,61,62,63,64,66,67,69,70,71,73,74,76,77,79,81,82,84,85,87,89,90,92,94,96,98,99,101,103,105,107,109,111,113,115,117,119,121,123,125,128,130,132,134,137,139,141,144,146,149,151,154,156,159,162,164,167,170,172,175,178,181,184,186,189,192,195,198,201,205,208,211,214,217,221,224,227,231,234,238,241,245,248,252,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,22,22,23,23,24,25,25,26,27,28,28,29,30,31,31,32,33,34,35,36,37,38,38,39,40,41,42,43,44,46,47,48,49,50,51,52,54,55,56,57,59,60,61,62,64,65,67,68,70,71,73,74,76,77,79,80,82,84,85,87,89,91,92,94,96,98,100,102,104,106,108,110,112,114,116,118,121,123,125,127,130,132,135,137,139,142,144,147,150,152,155,158,160,163,166,169,171,174,177,180,183,186,189,193,196,199,202,205,209,212,215,219,222,226,229,233,237,240,244,248,252,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,22,22,23,24,24,25,26,26,27,28,29,29,30,31,32,33,34,35,35,36,37,38,39,40,41,42,43,44,45,47,48,49,50,51,53,54,55,56,58,59,60,62,63,65,66,67,69,70,72,74,75,77,79,80,82,84,85,87,89,91,93,95,97,99,101,103,105,107,109,111,113,116,118,120,122,125,127,130,132,135,137,140,142,145,148,150,153,156,159,162,165,168,171,174,177,180,183,186,189,193,196,199,203,206,210,213,217,221,224,228,232,236,240,243,247,251,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,19,20,20,21,22,22,23,24,24,25,26,27,27,28,29,30,31,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,47,48,49,50,51,53,54,55,57,58,59,61,62,64,65,67,68,70,71,73,75,76,78,80,82,84,85,87,89,91,93,95,97,99,101,103,106,108,110,112,115,117,119,122,124,127,129,132,135,137,140,143,146,148,151,154,157,160,163,166,170,173,176,179,183,186,189,193,196,200,204,207,211,215,219,222,226,230,234,239,243,247,251,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,17,17,18,19,19,20,20,21,22,22,23,24,24,25,26,27,27,28,29,30,31,32,33,34,34,35,36,37,38,40,41,42,43,44,45,46,48,49,50,51,53,54,55,57,58,60,61,63,64,66,67,69,71,72,74,76,78,80,81,83,85,87,89,91,93,95,98,100,102,104,107,109,111,114,116,119,121,124,127,129,132,135,138,140,143,146,149,152,155,159,162,165,168,172,175,179,182,186,189,193,197,201,204,208,212,216,221,225,229,233,238,242,246,251,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,18,19,20,20,21,22,22,23,24,24,25,26,27,28,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,44,45,46,47,49,50,51,53,54,55,57,58,60,62,63,65,66,68,70,72,73,75,77,79,81,83,85,87,89,91,94,96,98,100,103,105,108,110,113,115,118,121,123,126,129,132,135,138,141,144,147,150,154,157,160,164,167,171,174,178,182,186,189,193,197,201,206,210,214,218,223,227,232,236,241,246,251,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,19,19,20,21,21,22,23,23,24,25,26,27,27,28,29,30,31,32,33,34,35,36,37,38,39,41,42,43,44,46,47,48,50,51,52,54,55,57,59,60,62,64,65,67,69,71,73,74,76,78,80,83,85,87,89,91,94,96,99,101,104,106,109,111,114,117,120,123,126,129,132,135,138,141,145,148,151,155,158,162,166,169,173,177,181,185,189,194,198,202,207,211,216,220,225,230,235,240,245,250,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15,16,16,17,17,18,19,19,20,21,22,22,23,24,25,25,26,27,28,29,30,31,32,33,34,35,36,37,39,40,41,42,44,45,46,48,49,51,52,54,55,57,59,60,62,64,66,68,69,71,73,76,78,80,82,84,87,89,91,94,96,99,102,104,107,110,113,116,119,122,125,128,131,135,138,142,145,149,153,156,160,164,168,172,176,181,185,189,194,199,203,208,213,218,223,228,233,239,244,250,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,12,12,12,13,13,14,15,15,16,16,17,17,18,19,19,20,21,22,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,38,39,40,41,43,44,46,47,49,50,52,53,55,57,58,60,62,64,66,68,70,72,74,77,79,81,84,86,89,91,94,97,99,102,105,108,111,114,118,121,124,128,131,135,138,142,146,150,154,158,162,166,171,175,180,185,189,194,199,204,210,215,220,226,232,237,243,249,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,5,6,6,6,7,7,7,7,8,8,8,9,9,10,10,10,11,11,12,12,13,13,14,14,15,15,16,17,17,18,19,19,20,21,22,23,23,24,25,26,27,28,29,30,31,33,34,35,36,37,39,40,42,43,45,46,48,49,51,53,55,56,58,60,62,64,66,69,71,73,75,78,80,83,86,88,91,94,97,100,103,106,109,113,116,120,123,127,131,135,139,143,147,151,155,160,165,169,174,179,184,189,195,200,206,212,217,223,229,236,242,249,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15,16,16,17,18,18,19,20,21,22,23,23,24,25,26,27,29,30,31,32,33,35,36,37,39,40,42,43,45,47,48,50,52,54,56,58,60,62,64,67,69,71,74,77,79,82,85,88,91,94,97,100,104,107,111,114,118,122,126,130,134,139,143,148,153,157,162,167,173,178,184,189,195,201,207,214,220,227,234,241,248,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11,12,12,13,13,14,14,15,16,16,17,18,19,20,21,21,22,23,24,25,27,28,29,30,31,33,34,35,37,38,40,42,43,45,47,49,51,53,55,57,60,62,64,67,69,72,75,78,81,84,87,90,94,97,101,104,108,112,116,121,125,129,134,139,144,149,154,160,165,171,177,183,189,196,203,210,217,224,232,239,247,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,9,9,10,10,11,11,12,12,13,14,14,15,16,16,17,18,19,20,21,22,23,24,25,26,28,29,30,32,33,35,36,38,40,42,43,45,47,49,52,54,56,59,61,64,67,70,73,76,79,82,86,89,93,97,101,105,110,114,119,124,129,134,139,145,150,156,163,169,175,182,189,197,204,212,220,229,237,246,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,4,5,5,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,14,15,15,16,17,18,19,20,21,22,24,25,26,27,29,30,32,34,35,37,39,41,43,45,48,50,52,55,58,61,64,67,70,73,77,81,84,88,93,97,101,106,111,116,122,127,133,139,146,152,159,166,174,181,189,198,206,216,225,235,245,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,10,10,11,12,12,13,14,15,16,17,18,19,20,21,23,24,25,27,29,30,32,34,36,38,40,43,45,48,50,53,56,59,63,66,70,74,78,82,87,92,97,102,107,113,119,126,132,139,147,155,163,171,180,189,199,209,220,231,243,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,9,9,10,11,11,12,13,14,15,16,17,18,20,21,23,24,26,28,30,32,34,36,39,41,44,47,51,54,58,61,66,70,74,79,85,90,96,102,109,116,123,131,140,148,158,168,178,189,201,214,227,241,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,9,9,10,11,11,12,13,14,15,16,17,18,20,21,23,24,26,28,30,32,34,36,39,41,44,47,51,54,58,61,66,70,74,79,85,90,96,102,109,116,123,131,140,148,158,168,178,189,201,214,227,241,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,9,9,10,11,11,12,13,14,15,16,17,18,20,21,23,24,26,28,30,32,34,36,39,41,44,47,51,54,58,61,66,70,74,79,85,90,96,102,109,116,123,131,140,148,158,168,178,189,201,214,227,241,255),
(0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,9,9,10,11,11,12,13,14,15,16,17,18,20,21,23,24,26,28,30,32,34,36,39,41,44,47,51,54,58,61,66,70,74,79,85,90,96,102,109,116,123,131,140,148,158,168,178,189,201,214,227,241,255));
type queue is array (0 to 255) of std_logic_vector (7 downto 0);
signal Q: queue;
signal flag : std_logic;
signal state : std_logic;
signal queue_index: std_logic_vector(7 DOWNTO 0);

begin

process(clk)
variable counter : integer range 0 to 255 :=0;
begin
  if(nrst = '1') then
    counter := 0;
	 flag <= '0';
	 state <= '0';
  elsif(rising_edge(clk)) then
	 Q(counter) <= input;
	 counter := counter+ 1;
	 if(counter = 256) then
	  counter := 0;
	  flag <= '1';
	end if;
	state <= not state;
  end if;
end process;
process(clk)
variable index : integer range 0 to 255 :=0;
begin
   if ( enable = '1') then
       output <= std_logic_vector(to_unsigned(lut(to_integer(unsigned(gamma)),to_integer(unsigned(Q(index)))),8));
		 index := index + 1;
		 queue_index <= Q(index);
		 if (index = 256) then
		     index := 0;
		 end if;
 end if;
end process;



end Behavioral;

